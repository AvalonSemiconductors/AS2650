// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire net91;
 wire clknet_leaf_0_wb_clk_i;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net92;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net93;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net94;
 wire net95;
 wire net80;
 wire net85;
 wire net81;
 wire net82;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net83;
 wire net84;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_3_0_wb_clk_i;
 wire clknet_opt_3_1_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4419_ (.I(net54),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4420_ (.I(\as2650.ins_reg[0] ),
    .Z(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4421_ (.I(_4001_),
    .Z(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4422_ (.I(_4002_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4423_ (.I(_4003_),
    .Z(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4424_ (.I(_4004_),
    .Z(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4425_ (.I(_4005_),
    .Z(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4426_ (.I(_4006_),
    .Z(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4427_ (.I(\as2650.psl[4] ),
    .Z(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4428_ (.I(_4008_),
    .Z(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4429_ (.I(_4009_),
    .Z(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4430_ (.I(_4010_),
    .Z(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4431_ (.I(_4011_),
    .Z(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4432_ (.I(_4012_),
    .Z(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4433_ (.I(_4013_),
    .Z(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4434_ (.I(_4014_),
    .ZN(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4435_ (.A1(\as2650.halted ),
    .A2(net10),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4436_ (.A1(_4015_),
    .A2(_4016_),
    .ZN(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4437_ (.I(_4001_),
    .Z(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4438_ (.I(\as2650.ins_reg[1] ),
    .Z(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4439_ (.A1(_4018_),
    .A2(_4019_),
    .ZN(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4440_ (.I(_4020_),
    .Z(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_4021_),
    .Z(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4442_ (.A1(_4017_),
    .A2(_4022_),
    .ZN(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4443_ (.I(_4023_),
    .Z(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4444_ (.I(\as2650.ins_reg[6] ),
    .Z(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4445_ (.I(_4025_),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4446_ (.I(_4026_),
    .Z(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4447_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(\as2650.cycle[5] ),
    .A4(\as2650.cycle[4] ),
    .ZN(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4448_ (.I(\as2650.cycle[3] ),
    .Z(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4449_ (.A1(_4029_),
    .A2(\as2650.cycle[2] ),
    .ZN(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4450_ (.A1(_4028_),
    .A2(_4030_),
    .ZN(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4451_ (.I(\as2650.cycle[1] ),
    .Z(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4452_ (.I(\as2650.cycle[0] ),
    .Z(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4453_ (.I(_4033_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4454_ (.I(_4034_),
    .Z(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(_4032_),
    .A2(_4035_),
    .ZN(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4456_ (.A1(_4031_),
    .A2(_4036_),
    .ZN(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4457_ (.I(_4037_),
    .Z(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4458_ (.I(\as2650.ins_reg[3] ),
    .Z(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4459_ (.I(_4039_),
    .ZN(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4460_ (.I(\as2650.ins_reg[4] ),
    .Z(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4461_ (.I(_4041_),
    .ZN(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4462_ (.I(_4042_),
    .Z(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4463_ (.A1(_4040_),
    .A2(_4043_),
    .ZN(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4464_ (.A1(_4027_),
    .A2(_4038_),
    .A3(_4044_),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4465_ (.I(\as2650.cycle[7] ),
    .Z(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4466_ (.I(_4046_),
    .ZN(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4467_ (.I(_4047_),
    .Z(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4468_ (.I(_4043_),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4469_ (.I(\as2650.cycle[5] ),
    .Z(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4470_ (.I(\as2650.cycle[6] ),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4471_ (.A1(_4051_),
    .A2(_4030_),
    .ZN(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4472_ (.I(\as2650.cycle[1] ),
    .ZN(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4473_ (.A1(_4053_),
    .A2(_4033_),
    .ZN(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4474_ (.A1(_4050_),
    .A2(\as2650.cycle[4] ),
    .A3(_4052_),
    .A4(_4054_),
    .ZN(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4475_ (.I(_4055_),
    .Z(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4476_ (.I(\as2650.idx_ctrl[1] ),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4477_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4478_ (.A1(_4057_),
    .A2(_4058_),
    .ZN(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4479_ (.I(_4059_),
    .Z(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4480_ (.A1(_4048_),
    .A2(_4049_),
    .A3(_4056_),
    .A4(_4060_),
    .ZN(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4481_ (.I(\as2650.ins_reg[2] ),
    .Z(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4482_ (.I(_4062_),
    .Z(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4483_ (.I(\as2650.ins_reg[5] ),
    .Z(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4484_ (.I(_4064_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4485_ (.I(_4065_),
    .ZN(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4486_ (.I(_4041_),
    .Z(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4487_ (.A1(_4066_),
    .A2(_4067_),
    .ZN(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4488_ (.I(\as2650.ins_reg[7] ),
    .Z(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4489_ (.I(_4069_),
    .ZN(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4490_ (.A1(_4026_),
    .A2(_4070_),
    .ZN(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4491_ (.A1(_4063_),
    .A2(_4068_),
    .A3(_4071_),
    .Z(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4492_ (.I(_4063_),
    .Z(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4493_ (.A1(_4025_),
    .A2(\as2650.ins_reg[7] ),
    .ZN(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4494_ (.A1(_4064_),
    .A2(_4074_),
    .ZN(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4495_ (.A1(_4041_),
    .A2(_4075_),
    .ZN(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4496_ (.I(_4076_),
    .Z(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4497_ (.A1(_4073_),
    .A2(_4077_),
    .Z(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4498_ (.A1(_4072_),
    .A2(_4078_),
    .ZN(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4499_ (.I(_4039_),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4500_ (.A1(_4053_),
    .A2(_4031_),
    .ZN(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4501_ (.A1(_4034_),
    .A2(_4081_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4502_ (.I(_4082_),
    .Z(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4503_ (.A1(_4080_),
    .A2(_4083_),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4504_ (.A1(_4079_),
    .A2(_4084_),
    .ZN(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4505_ (.A1(_4045_),
    .A2(_4061_),
    .A3(_4085_),
    .ZN(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(_4067_),
    .Z(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4507_ (.I(_4087_),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4508_ (.I(_4088_),
    .Z(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4509_ (.I(_4046_),
    .Z(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4510_ (.A1(_4090_),
    .A2(_4055_),
    .ZN(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4511_ (.I(_4091_),
    .Z(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4512_ (.I(\as2650.addr_buff[7] ),
    .Z(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4513_ (.I(\as2650.addr_buff[6] ),
    .Z(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4514_ (.I(\as2650.addr_buff[5] ),
    .Z(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4515_ (.A1(_4094_),
    .A2(_4095_),
    .ZN(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4516_ (.A1(_4093_),
    .A2(_4096_),
    .Z(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4517_ (.A1(_4089_),
    .A2(_4092_),
    .A3(_4097_),
    .ZN(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4518_ (.A1(_4065_),
    .A2(_4041_),
    .ZN(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4519_ (.A1(_4062_),
    .A2(_4099_),
    .ZN(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4520_ (.A1(_4070_),
    .A2(_4100_),
    .ZN(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4521_ (.I(_4028_),
    .Z(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4522_ (.A1(\as2650.cycle[1] ),
    .A2(\as2650.cycle[0] ),
    .Z(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4523_ (.A1(_4102_),
    .A2(_4030_),
    .A3(_4103_),
    .ZN(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4524_ (.I(_4104_),
    .Z(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4525_ (.A1(_4039_),
    .A2(_4101_),
    .A3(_4105_),
    .ZN(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4526_ (.A1(_4086_),
    .A2(_4098_),
    .A3(_4106_),
    .Z(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4527_ (.I(_4083_),
    .Z(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4528_ (.I(_4108_),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4529_ (.I(_4016_),
    .Z(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4530_ (.A1(_4014_),
    .A2(_4022_),
    .ZN(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4531_ (.A1(_4110_),
    .A2(_4111_),
    .ZN(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4532_ (.A1(_4062_),
    .A2(\as2650.ins_reg[3] ),
    .ZN(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4533_ (.I(_4113_),
    .Z(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4534_ (.I(_4114_),
    .Z(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4535_ (.A1(_4043_),
    .A2(_4115_),
    .A3(_4075_),
    .ZN(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4536_ (.A1(_4109_),
    .A2(_4112_),
    .A3(_4116_),
    .ZN(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4537_ (.I(_4033_),
    .Z(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4538_ (.I(\as2650.cycle[1] ),
    .Z(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4539_ (.I(\as2650.cycle[3] ),
    .ZN(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4540_ (.I(\as2650.cycle[2] ),
    .Z(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4541_ (.A1(_4120_),
    .A2(_4121_),
    .A3(_4028_),
    .ZN(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4542_ (.A1(_4119_),
    .A2(_4122_),
    .Z(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4543_ (.A1(_4118_),
    .A2(_4123_),
    .ZN(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4544_ (.I(_4124_),
    .Z(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4545_ (.A1(_4064_),
    .A2(_4026_),
    .A3(_4069_),
    .ZN(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4546_ (.I(_4126_),
    .Z(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4547_ (.I(_4087_),
    .Z(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4548_ (.I(_4115_),
    .Z(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4549_ (.A1(_4128_),
    .A2(_4129_),
    .ZN(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4550_ (.I(_4022_),
    .Z(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4551_ (.A1(_4131_),
    .A2(_4059_),
    .ZN(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4552_ (.A1(_4125_),
    .A2(_4127_),
    .A3(_4130_),
    .A4(_4132_),
    .ZN(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4553_ (.A1(_4017_),
    .A2(_4133_),
    .ZN(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_4134_),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4555_ (.A1(_4024_),
    .A2(_4107_),
    .B(_4117_),
    .C(_4135_),
    .ZN(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4556_ (.A1(_4007_),
    .A2(_4136_),
    .Z(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4557_ (.I(_4137_),
    .Z(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4558_ (.I(_4135_),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4559_ (.I(_4065_),
    .Z(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4560_ (.I(_4140_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4561_ (.I(_4141_),
    .Z(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4562_ (.I(_4069_),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4563_ (.A1(_4026_),
    .A2(_4143_),
    .ZN(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4564_ (.I(_4144_),
    .Z(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4565_ (.A1(_4142_),
    .A2(_4145_),
    .ZN(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4566_ (.I(_4146_),
    .Z(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4567_ (.I(\as2650.r0[0] ),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4568_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_4009_),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4569_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123_2[1][0] ),
    .S(_4010_),
    .Z(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4570_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_4009_),
    .Z(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4571_ (.I0(_4148_),
    .I1(_4149_),
    .I2(_4150_),
    .I3(_4151_),
    .S0(_4018_),
    .S1(_4019_),
    .Z(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4572_ (.I(_4152_),
    .Z(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4573_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4574_ (.A1(\as2650.holding_reg[0] ),
    .A2(_4154_),
    .Z(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4575_ (.A1(_4113_),
    .A2(_4153_),
    .B(_4155_),
    .ZN(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4576_ (.I0(\as2650.holding_reg[0] ),
    .I1(_4153_),
    .S(_4154_),
    .Z(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4577_ (.A1(_4156_),
    .A2(_4157_),
    .Z(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4578_ (.I(_4158_),
    .Z(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4579_ (.I(_4152_),
    .Z(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_4160_),
    .Z(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4581_ (.A1(\as2650.holding_reg[0] ),
    .A2(_4161_),
    .ZN(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4582_ (.I(_4140_),
    .Z(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4583_ (.I(_4071_),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4584_ (.A1(_4163_),
    .A2(_4164_),
    .ZN(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4585_ (.I(_4025_),
    .ZN(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4586_ (.A1(_4166_),
    .A2(_4143_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4587_ (.I(_4167_),
    .Z(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4588_ (.I(_4157_),
    .Z(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4589_ (.A1(_4027_),
    .A2(_4070_),
    .ZN(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4590_ (.I(_4170_),
    .Z(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4591_ (.A1(_4141_),
    .A2(_4171_),
    .ZN(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4592_ (.I(\as2650.carry ),
    .ZN(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4593_ (.A1(\as2650.psl[3] ),
    .A2(_4173_),
    .ZN(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4594_ (.I(_4174_),
    .ZN(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4595_ (.A1(_4175_),
    .A2(_4158_),
    .Z(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(\as2650.psl[3] ),
    .A2(\as2650.carry ),
    .ZN(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4597_ (.I(_4066_),
    .Z(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4598_ (.A1(_4178_),
    .A2(_4170_),
    .ZN(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4599_ (.A1(_4177_),
    .A2(_4158_),
    .B(_4179_),
    .ZN(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4600_ (.A1(_4177_),
    .A2(_4159_),
    .B(_4180_),
    .ZN(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4601_ (.A1(_4171_),
    .A2(_4156_),
    .B1(_4172_),
    .B2(_4176_),
    .C(_4181_),
    .ZN(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4602_ (.A1(_4168_),
    .A2(_4169_),
    .B(_4165_),
    .C(_4182_),
    .ZN(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4603_ (.A1(_4162_),
    .A2(_4165_),
    .B(_4183_),
    .ZN(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4604_ (.A1(_4147_),
    .A2(_4184_),
    .ZN(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4605_ (.A1(_4147_),
    .A2(_4159_),
    .B(_4185_),
    .ZN(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4606_ (.I(_4148_),
    .Z(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4607_ (.I(_4187_),
    .Z(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4608_ (.I(_4188_),
    .Z(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4609_ (.I(_4154_),
    .Z(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4610_ (.I(_4190_),
    .Z(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4611_ (.I(_4191_),
    .Z(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_4192_),
    .Z(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4613_ (.I(_4075_),
    .Z(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(_4043_),
    .A2(_4194_),
    .ZN(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4615_ (.A1(_4193_),
    .A2(_4195_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4616_ (.A1(_4082_),
    .A2(_4112_),
    .ZN(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4617_ (.A1(_4196_),
    .A2(_4197_),
    .ZN(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4618_ (.I(_4198_),
    .Z(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4619_ (.I(_4199_),
    .Z(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4620_ (.I(_4199_),
    .Z(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4621_ (.A1(_4192_),
    .A2(_4077_),
    .ZN(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4622_ (.A1(_4202_),
    .A2(_4197_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4623_ (.I(_4203_),
    .Z(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4624_ (.I(_4204_),
    .Z(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4625_ (.I(\as2650.psl[3] ),
    .Z(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4626_ (.I(_4206_),
    .ZN(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4627_ (.I(\as2650.r0[7] ),
    .Z(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4628_ (.I(_4208_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4629_ (.I(_4209_),
    .Z(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4630_ (.A1(_4210_),
    .A2(_4022_),
    .ZN(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4631_ (.A1(_4001_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4632_ (.I(_4212_),
    .Z(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4633_ (.I(_4213_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4634_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_4013_),
    .Z(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4635_ (.A1(_4214_),
    .A2(_4215_),
    .ZN(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4636_ (.A1(\as2650.ins_reg[0] ),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4637_ (.I(_4217_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4638_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_4003_),
    .S1(_4014_),
    .Z(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4639_ (.A1(_4218_),
    .A2(_4219_),
    .ZN(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4640_ (.A1(_4211_),
    .A2(_4216_),
    .A3(_4220_),
    .Z(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4641_ (.I(_4221_),
    .Z(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4642_ (.I(_4222_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4643_ (.A1(_4207_),
    .A2(_4223_),
    .B(_4175_),
    .ZN(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4644_ (.A1(_4080_),
    .A2(_4072_),
    .ZN(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4645_ (.A1(_4225_),
    .A2(_4197_),
    .ZN(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4646_ (.I(_4226_),
    .Z(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(_4227_),
    .Z(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4648_ (.I(\as2650.r0[1] ),
    .Z(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4649_ (.I(_4229_),
    .ZN(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4650_ (.A1(_4001_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4651_ (.A1(_4230_),
    .A2(_4231_),
    .ZN(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4652_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_4010_),
    .Z(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4653_ (.A1(_4212_),
    .A2(_4233_),
    .Z(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4654_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_4010_),
    .Z(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4655_ (.A1(_4217_),
    .A2(_4235_),
    .Z(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4656_ (.A1(_4232_),
    .A2(_4234_),
    .A3(_4236_),
    .ZN(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4657_ (.I(_4237_),
    .Z(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4658_ (.I(_4238_),
    .Z(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4659_ (.I(_4203_),
    .Z(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4660_ (.I(net5),
    .Z(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4661_ (.I(_4241_),
    .Z(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4662_ (.I(_4242_),
    .Z(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4663_ (.A1(_4023_),
    .A2(_4106_),
    .ZN(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4664_ (.I(_4244_),
    .Z(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4665_ (.I(_4245_),
    .Z(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4666_ (.I(_4244_),
    .Z(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4667_ (.A1(\as2650.ins_reg[4] ),
    .A2(_4025_),
    .A3(\as2650.ins_reg[7] ),
    .ZN(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4668_ (.I(_4161_),
    .Z(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4669_ (.A1(_4248_),
    .A2(_4249_),
    .Z(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4670_ (.A1(_4247_),
    .A2(_4250_),
    .ZN(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4671_ (.I(_4226_),
    .Z(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4672_ (.A1(_4243_),
    .A2(_4246_),
    .B(_4251_),
    .C(_4252_),
    .ZN(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4673_ (.A1(_4228_),
    .A2(_4239_),
    .B(_4240_),
    .C(_4253_),
    .ZN(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4674_ (.A1(_4205_),
    .A2(_4224_),
    .B(_4254_),
    .ZN(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4675_ (.A1(_4201_),
    .A2(_4255_),
    .ZN(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4676_ (.A1(_4024_),
    .A2(_4098_),
    .ZN(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4677_ (.I(_4257_),
    .Z(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4678_ (.A1(_4189_),
    .A2(_4200_),
    .B(_4256_),
    .C(_4258_),
    .ZN(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4679_ (.I(_4088_),
    .Z(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4680_ (.A1(_4260_),
    .A2(_4092_),
    .ZN(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4681_ (.A1(_4093_),
    .A2(_4096_),
    .ZN(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4682_ (.A1(_4261_),
    .A2(_4262_),
    .ZN(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4683_ (.A1(_4112_),
    .A2(_4263_),
    .ZN(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4684_ (.I(_4153_),
    .Z(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4685_ (.I(\as2650.addr_buff[5] ),
    .ZN(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4686_ (.A1(\as2650.addr_buff[6] ),
    .A2(_4266_),
    .ZN(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4687_ (.I(\as2650.addr_buff[6] ),
    .ZN(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4688_ (.A1(_4268_),
    .A2(\as2650.addr_buff[5] ),
    .ZN(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4689_ (.A1(_4267_),
    .A2(_4269_),
    .ZN(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4690_ (.A1(_4265_),
    .A2(_4270_),
    .ZN(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4691_ (.I(_4271_),
    .Z(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4692_ (.A1(_4112_),
    .A2(_4061_),
    .ZN(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4693_ (.A1(_4264_),
    .A2(_4272_),
    .B(_4273_),
    .ZN(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4694_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_4058_),
    .ZN(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4695_ (.A1(_4057_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4696_ (.A1(_4275_),
    .A2(_4276_),
    .ZN(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4697_ (.A1(_4265_),
    .A2(_4277_),
    .Z(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4698_ (.I(_4278_),
    .Z(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4699_ (.I(_4273_),
    .Z(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4700_ (.I(_4135_),
    .Z(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4701_ (.A1(_4259_),
    .A2(_4274_),
    .B1(_4279_),
    .B2(_4280_),
    .C(_4281_),
    .ZN(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4702_ (.A1(_4139_),
    .A2(_4186_),
    .B(_4282_),
    .ZN(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4703_ (.I(net10),
    .ZN(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4704_ (.I(_4284_),
    .Z(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4705_ (.I(_4014_),
    .Z(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4706_ (.I(\as2650.halted ),
    .ZN(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4707_ (.A1(_4287_),
    .A2(_4284_),
    .ZN(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4708_ (.A1(_4286_),
    .A2(_4288_),
    .ZN(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4709_ (.I(_4289_),
    .Z(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4710_ (.I(_4037_),
    .Z(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4711_ (.I(_4291_),
    .Z(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4712_ (.I(_4292_),
    .Z(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4713_ (.I(_4293_),
    .Z(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4714_ (.I(_4115_),
    .Z(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4715_ (.A1(_4131_),
    .A2(_4295_),
    .ZN(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4716_ (.A1(_4166_),
    .A2(_4069_),
    .ZN(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4717_ (.I(_4297_),
    .Z(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4718_ (.I(_4298_),
    .Z(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4719_ (.I(_4068_),
    .Z(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4720_ (.A1(_4296_),
    .A2(_4299_),
    .A3(_4300_),
    .ZN(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4721_ (.A1(_4290_),
    .A2(_4294_),
    .A3(_4301_),
    .ZN(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4722_ (.A1(_4285_),
    .A2(_4302_),
    .A3(_4137_),
    .Z(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4723_ (.I(_4303_),
    .Z(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4724_ (.A1(\as2650.r123[1][0] ),
    .A2(_4304_),
    .ZN(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4725_ (.I(_4189_),
    .Z(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4726_ (.I(_4291_),
    .Z(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4727_ (.I(_4307_),
    .Z(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4728_ (.A1(_4289_),
    .A2(_4308_),
    .ZN(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4729_ (.I(_4231_),
    .Z(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4730_ (.A1(_4310_),
    .A2(_4192_),
    .ZN(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4731_ (.A1(_4297_),
    .A2(_4300_),
    .ZN(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4732_ (.A1(_4311_),
    .A2(_4312_),
    .ZN(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4733_ (.I(_4313_),
    .Z(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4734_ (.A1(_4309_),
    .A2(_4314_),
    .ZN(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4735_ (.I(_4315_),
    .Z(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4736_ (.I(_4316_),
    .Z(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4737_ (.I(_4149_),
    .Z(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4738_ (.I(_4318_),
    .Z(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4739_ (.I(_4319_),
    .Z(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4740_ (.I(_4320_),
    .Z(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4741_ (.I(_4321_),
    .Z(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4742_ (.A1(_4306_),
    .A2(_4317_),
    .A3(_4322_),
    .ZN(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4743_ (.A1(_4138_),
    .A2(_4283_),
    .B(_4305_),
    .C(_4323_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4744_ (.I(_4137_),
    .Z(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4745_ (.A1(_4163_),
    .A2(_4145_),
    .Z(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4746_ (.I(\as2650.holding_reg[1] ),
    .Z(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4747_ (.A1(_4326_),
    .A2(_4113_),
    .ZN(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4748_ (.A1(_4114_),
    .A2(_4238_),
    .B(_4327_),
    .ZN(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4749_ (.I(_4328_),
    .Z(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4750_ (.A1(_4325_),
    .A2(_4329_),
    .ZN(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4751_ (.A1(_4178_),
    .A2(_4167_),
    .ZN(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4752_ (.A1(_4232_),
    .A2(_4234_),
    .A3(_4236_),
    .Z(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4753_ (.A1(\as2650.holding_reg[1] ),
    .A2(_4332_),
    .Z(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4754_ (.I(_4333_),
    .Z(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4755_ (.A1(_4178_),
    .A2(_4298_),
    .ZN(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4756_ (.A1(\as2650.holding_reg[1] ),
    .A2(_4332_),
    .ZN(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4757_ (.A1(_4334_),
    .A2(_4336_),
    .ZN(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4758_ (.A1(_4156_),
    .A2(_4157_),
    .ZN(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4759_ (.A1(_4162_),
    .A2(_4169_),
    .ZN(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4760_ (.A1(_4175_),
    .A2(_4338_),
    .B(_4339_),
    .ZN(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4761_ (.A1(_4337_),
    .A2(_4340_),
    .Z(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4762_ (.A1(_4335_),
    .A2(_4341_),
    .ZN(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4763_ (.A1(_4065_),
    .A2(_4298_),
    .ZN(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4764_ (.A1(_4333_),
    .A2(_4336_),
    .Z(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4765_ (.A1(_4177_),
    .A2(_4158_),
    .B(_4162_),
    .ZN(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4766_ (.A1(_4344_),
    .A2(_4345_),
    .Z(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4767_ (.A1(_4343_),
    .A2(_4346_),
    .ZN(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4768_ (.A1(_4140_),
    .A2(_4168_),
    .ZN(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4769_ (.A1(_4326_),
    .A2(_4191_),
    .ZN(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4770_ (.A1(_4192_),
    .A2(_4239_),
    .B(_4349_),
    .C(_4298_),
    .ZN(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4771_ (.A1(_4342_),
    .A2(_4347_),
    .A3(_4348_),
    .A4(_4350_),
    .Z(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4772_ (.A1(_4141_),
    .A2(_4336_),
    .B(_4164_),
    .ZN(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4773_ (.A1(_4331_),
    .A2(_4334_),
    .B1(_4351_),
    .B2(_4352_),
    .ZN(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4774_ (.A1(_4330_),
    .A2(_4353_),
    .ZN(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4775_ (.I(_4354_),
    .ZN(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4776_ (.A1(_4057_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4777_ (.A1(_4161_),
    .A2(_4356_),
    .B(_4276_),
    .ZN(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4778_ (.A1(_4161_),
    .A2(_4237_),
    .A3(_4357_),
    .Z(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4779_ (.I(_4358_),
    .Z(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4780_ (.A1(_4280_),
    .A2(_4359_),
    .ZN(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4781_ (.I(_4088_),
    .Z(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4782_ (.I(_4361_),
    .Z(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4783_ (.A1(_4048_),
    .A2(_4055_),
    .ZN(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4784_ (.I(_4363_),
    .Z(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4785_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4786_ (.A1(_4362_),
    .A2(_4364_),
    .A3(_4365_),
    .ZN(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4787_ (.A1(_4024_),
    .A2(_4366_),
    .ZN(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4788_ (.I(_4367_),
    .Z(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4789_ (.I(_4257_),
    .Z(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4790_ (.I(_4369_),
    .Z(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4791_ (.A1(_4268_),
    .A2(\as2650.addr_buff[5] ),
    .ZN(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4792_ (.A1(_4160_),
    .A2(_4371_),
    .B(_4269_),
    .ZN(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4793_ (.A1(_4160_),
    .A2(_4332_),
    .A3(_4372_),
    .Z(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4794_ (.I(_4373_),
    .Z(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4795_ (.I(_4229_),
    .Z(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4796_ (.I(_4375_),
    .Z(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4797_ (.I(_4376_),
    .Z(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4798_ (.I(_4198_),
    .Z(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4799_ (.I(_4249_),
    .Z(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4800_ (.I(_4203_),
    .Z(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(\as2650.r0[2] ),
    .Z(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4802_ (.I(_4381_),
    .Z(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4803_ (.A1(_4382_),
    .A2(_4020_),
    .ZN(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4804_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_4011_),
    .Z(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4805_ (.A1(_4212_),
    .A2(_4384_),
    .ZN(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4806_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_4018_),
    .S1(_4011_),
    .Z(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4807_ (.A1(_4217_),
    .A2(_4386_),
    .ZN(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4808_ (.A1(_4383_),
    .A2(_4385_),
    .A3(_4387_),
    .ZN(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4809_ (.I(_4388_),
    .Z(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4810_ (.I(_4389_),
    .Z(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4811_ (.I(net6),
    .Z(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4812_ (.I(_4391_),
    .Z(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4813_ (.I(_4392_),
    .Z(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4814_ (.A1(_4064_),
    .A2(_4248_),
    .ZN(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4815_ (.A1(_4394_),
    .A2(_4249_),
    .ZN(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4816_ (.A1(\as2650.ins_reg[5] ),
    .A2(\as2650.ins_reg[6] ),
    .A3(\as2650.ins_reg[7] ),
    .Z(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4817_ (.A1(\as2650.ins_reg[4] ),
    .A2(_4396_),
    .ZN(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4818_ (.A1(_4265_),
    .A2(_4397_),
    .Z(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4819_ (.A1(_4395_),
    .A2(_4398_),
    .ZN(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4820_ (.A1(_4238_),
    .A2(_4399_),
    .Z(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4821_ (.A1(_4244_),
    .A2(_4400_),
    .ZN(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4822_ (.A1(_4393_),
    .A2(_4245_),
    .B(_4401_),
    .ZN(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4823_ (.A1(_4227_),
    .A2(_4402_),
    .ZN(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4824_ (.A1(_4252_),
    .A2(_4390_),
    .B(_4403_),
    .ZN(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4825_ (.A1(_4240_),
    .A2(_4404_),
    .ZN(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4826_ (.A1(_4379_),
    .A2(_4380_),
    .B(_4405_),
    .ZN(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4827_ (.A1(_4378_),
    .A2(_4406_),
    .ZN(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4828_ (.A1(_4377_),
    .A2(_4201_),
    .B(_4369_),
    .C(_4407_),
    .ZN(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4829_ (.A1(_4370_),
    .A2(_4374_),
    .B(_4408_),
    .ZN(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4830_ (.A1(_4368_),
    .A2(_4409_),
    .ZN(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4831_ (.A1(_4360_),
    .A2(_4410_),
    .B(_4281_),
    .ZN(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4832_ (.A1(_4139_),
    .A2(_4355_),
    .B(_4411_),
    .ZN(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(_4303_),
    .Z(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4834_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_4008_),
    .Z(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4835_ (.I(_4414_),
    .Z(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4836_ (.I(_4415_),
    .Z(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4837_ (.I(_4416_),
    .Z(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4838_ (.A1(_4376_),
    .A2(_4188_),
    .A3(_4321_),
    .A4(_4417_),
    .ZN(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4839_ (.I(_4418_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4840_ (.A1(_4377_),
    .A2(_4322_),
    .B1(_4417_),
    .B2(_4189_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4841_ (.A1(_0284_),
    .A2(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4842_ (.I(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4843_ (.I(_4315_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4844_ (.A1(\as2650.r123[1][1] ),
    .A2(_4413_),
    .B1(_0287_),
    .B2(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4845_ (.A1(_4324_),
    .A2(_4412_),
    .B(_0289_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4846_ (.I(_4125_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4847_ (.A1(_0290_),
    .A2(_4127_),
    .A3(_4130_),
    .A4(_4132_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4848_ (.A1(_4289_),
    .A2(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4849_ (.I(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4850_ (.I(_4388_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4851_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0294_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4852_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0294_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4853_ (.A1(_0295_),
    .A2(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4854_ (.I(_0297_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4855_ (.I(_4165_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4856_ (.A1(_4383_),
    .A2(_4385_),
    .A3(_4387_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4857_ (.I(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(\as2650.holding_reg[2] ),
    .A2(_4190_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4859_ (.A1(_4190_),
    .A2(_0301_),
    .B(_0302_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4860_ (.I(_4332_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4861_ (.A1(_4326_),
    .A2(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4862_ (.A1(_4328_),
    .A2(_0305_),
    .B1(_4344_),
    .B2(_4340_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4863_ (.A1(_0297_),
    .A2(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4864_ (.A1(_4337_),
    .A2(_4345_),
    .B(_4334_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4865_ (.A1(_0298_),
    .A2(_0308_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4866_ (.A1(_4335_),
    .A2(_0307_),
    .B1(_0309_),
    .B2(_4343_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4867_ (.A1(_4171_),
    .A2(_0303_),
    .B(_0310_),
    .C(_4348_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4868_ (.I(_4168_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4869_ (.A1(_4178_),
    .A2(_0296_),
    .B(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4870_ (.A1(_0299_),
    .A2(_0295_),
    .B1(_0311_),
    .B2(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4871_ (.I0(_0298_),
    .I1(_0314_),
    .S(_4146_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4872_ (.I(_0315_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4873_ (.I(_4367_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4874_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_4058_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4875_ (.A1(_4160_),
    .A2(_4232_),
    .A3(_4234_),
    .A4(_4236_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4876_ (.A1(_0319_),
    .A2(_4388_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4877_ (.A1(_0318_),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4878_ (.A1(_4356_),
    .A2(_0318_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _4879_ (.A1(_4232_),
    .A2(_4234_),
    .A3(_4236_),
    .B(_4153_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4880_ (.I(_0300_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4881_ (.A1(_0323_),
    .A2(_0324_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4882_ (.A1(_0322_),
    .A2(_4389_),
    .B1(_0325_),
    .B2(_4356_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4883_ (.A1(_0321_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4884_ (.A1(\as2650.addr_buff[6] ),
    .A2(_4266_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4885_ (.A1(_4270_),
    .A2(_0301_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4886_ (.A1(_0328_),
    .A2(_0320_),
    .B1(_0325_),
    .B2(_4371_),
    .C(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4887_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4888_ (.I(_4382_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4889_ (.I(_0332_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4890_ (.I(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4891_ (.I(\as2650.r0[3] ),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4892_ (.I(_0335_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4893_ (.I(_0336_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4894_ (.A1(_0337_),
    .A2(_4020_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4895_ (.I(_4011_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4896_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4897_ (.A1(_4213_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4898_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_4018_),
    .S1(_0339_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4899_ (.A1(_4218_),
    .A2(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4900_ (.A1(_0338_),
    .A2(_0341_),
    .A3(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4901_ (.I(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4902_ (.I(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4903_ (.I(net7),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4904_ (.I(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4905_ (.I(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4906_ (.A1(_4143_),
    .A2(_4099_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4907_ (.A1(_4063_),
    .A2(_4104_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4908_ (.A1(_0350_),
    .A2(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4909_ (.A1(_4039_),
    .A2(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4910_ (.A1(_4024_),
    .A2(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4911_ (.I(_0324_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4912_ (.I0(_4395_),
    .I1(_4398_),
    .S(_4238_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4913_ (.A1(_0355_),
    .A2(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(_0354_),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4915_ (.A1(_0349_),
    .A2(_0354_),
    .B(_0358_),
    .C(_4226_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4916_ (.A1(_4252_),
    .A2(_0346_),
    .B(_0359_),
    .C(_4203_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4917_ (.A1(_4240_),
    .A2(_4239_),
    .B(_0360_),
    .C(_4198_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4918_ (.A1(_0334_),
    .A2(_4199_),
    .B(_4257_),
    .C(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4919_ (.A1(_4258_),
    .A2(_0331_),
    .B(_0362_),
    .C(_4367_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4920_ (.A1(_0317_),
    .A2(_0327_),
    .B(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4921_ (.A1(_0292_),
    .A2(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4922_ (.A1(_0293_),
    .A2(_0316_),
    .B(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4923_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(_4008_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4924_ (.I(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4925_ (.I(_0368_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4926_ (.I(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4927_ (.A1(_4187_),
    .A2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4928_ (.I(_4415_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4929_ (.I(_4375_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4930_ (.A1(_0333_),
    .A2(_4320_),
    .B1(_0372_),
    .B2(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4931_ (.A1(_0332_),
    .A2(_0373_),
    .A3(_4320_),
    .A4(_0372_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4932_ (.A1(_0371_),
    .A2(_0374_),
    .A3(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4933_ (.A1(_0374_),
    .A2(_0375_),
    .B(_0371_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4934_ (.A1(_0284_),
    .A2(_0376_),
    .A3(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4935_ (.A1(_0376_),
    .A2(_0377_),
    .B(_0284_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4936_ (.A1(_0378_),
    .A2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4937_ (.A1(\as2650.r123[1][2] ),
    .A2(_4413_),
    .B1(_0380_),
    .B2(_4316_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4938_ (.A1(_4324_),
    .A2(_0366_),
    .B(_0381_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4939_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0344_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4940_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0345_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4941_ (.A1(_0382_),
    .A2(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4942_ (.I(_4335_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4943_ (.A1(_0382_),
    .A2(_0383_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4944_ (.I(\as2650.holding_reg[2] ),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4945_ (.A1(_0387_),
    .A2(_0294_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4946_ (.A1(_0297_),
    .A2(_0306_),
    .B1(_0303_),
    .B2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4947_ (.A1(_0386_),
    .A2(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4948_ (.A1(_0385_),
    .A2(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4949_ (.A1(_0387_),
    .A2(_4389_),
    .B1(_4337_),
    .B2(_4345_),
    .C(_4334_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4950_ (.A1(_0388_),
    .A2(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4951_ (.A1(_0384_),
    .A2(_0393_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4952_ (.I(\as2650.holding_reg[3] ),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4953_ (.I(_4115_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4954_ (.I(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4955_ (.A1(_0338_),
    .A2(_0341_),
    .A3(_0343_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4956_ (.I(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4957_ (.I(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4958_ (.A1(_4129_),
    .A2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4959_ (.A1(_0395_),
    .A2(_0397_),
    .B(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4960_ (.I(_4299_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4961_ (.A1(_4343_),
    .A2(_0394_),
    .B1(_0402_),
    .B2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4962_ (.I(_4142_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4963_ (.A1(_4190_),
    .A2(_0399_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4964_ (.A1(_0395_),
    .A2(_4191_),
    .B(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4965_ (.A1(_0405_),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4966_ (.A1(_0391_),
    .A2(_0404_),
    .B1(_0408_),
    .B2(_0312_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4967_ (.I(_4331_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4968_ (.A1(_0410_),
    .A2(_0382_),
    .B(_4146_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4969_ (.A1(_4147_),
    .A2(_0384_),
    .B1(_0409_),
    .B2(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4970_ (.I(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4971_ (.I(_0337_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4972_ (.I(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4973_ (.I(\as2650.r0[4] ),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4974_ (.I(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4975_ (.I(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4976_ (.A1(_0418_),
    .A2(_4021_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4977_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_0339_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4978_ (.A1(_4213_),
    .A2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4979_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_4002_),
    .S1(_0339_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4980_ (.A1(_4218_),
    .A2(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _4981_ (.A1(_0419_),
    .A2(_0421_),
    .A3(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4982_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4983_ (.I(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4984_ (.I(_0426_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4985_ (.I(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4986_ (.I(net8),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4987_ (.I(_0429_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4988_ (.I(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4989_ (.I(_4226_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4990_ (.A1(_4076_),
    .A2(_0323_),
    .A3(_0301_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4991_ (.A1(_0304_),
    .A2(_4398_),
    .A3(_0294_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4992_ (.A1(_0433_),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4993_ (.A1(_0346_),
    .A2(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4994_ (.A1(_4247_),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4995_ (.A1(_0431_),
    .A2(_4246_),
    .B(_0432_),
    .C(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4996_ (.A1(_4228_),
    .A2(_0428_),
    .B(_0438_),
    .C(_4380_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4997_ (.A1(_4205_),
    .A2(_4390_),
    .B(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4998_ (.A1(_4201_),
    .A2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4999_ (.A1(_0415_),
    .A2(_4200_),
    .B(_4370_),
    .C(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5000_ (.I(_4270_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5001_ (.A1(_0319_),
    .A2(_0324_),
    .A3(_0398_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5002_ (.A1(_0319_),
    .A2(_0301_),
    .B(_0399_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5003_ (.A1(_0444_),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5004_ (.I(_4269_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5005_ (.A1(_4265_),
    .A2(_0304_),
    .A3(_4388_),
    .A4(_0344_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5006_ (.A1(_0323_),
    .A2(_0324_),
    .B(_0399_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5007_ (.A1(_0448_),
    .A2(_0449_),
    .B(_4371_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5008_ (.A1(_0443_),
    .A2(_0400_),
    .B1(_0446_),
    .B2(_0447_),
    .C(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5009_ (.I(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5010_ (.A1(_4264_),
    .A2(_0452_),
    .B(_4273_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5011_ (.I(_4277_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5012_ (.I(_4276_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5013_ (.A1(_0448_),
    .A2(_0449_),
    .B(_4356_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5014_ (.A1(_0454_),
    .A2(_0400_),
    .B1(_0446_),
    .B2(_0455_),
    .C(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5015_ (.I(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5016_ (.A1(_0317_),
    .A2(_0458_),
    .B(_0292_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5017_ (.A1(_0442_),
    .A2(_0453_),
    .B(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5018_ (.A1(_4139_),
    .A2(_0413_),
    .B(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5019_ (.I(_4302_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5020_ (.A1(_0284_),
    .A2(_0376_),
    .A3(_0377_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5021_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(_4008_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5022_ (.I(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5023_ (.I(_0465_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5024_ (.I(_0466_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5025_ (.A1(_4375_),
    .A2(_4187_),
    .A3(_0370_),
    .A4(_0467_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5026_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5027_ (.I(_0467_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5028_ (.A1(_0373_),
    .A2(_0370_),
    .B1(_0470_),
    .B2(_4187_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5029_ (.A1(_0414_),
    .A2(_4319_),
    .B1(_4416_),
    .B2(_0332_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5030_ (.A1(_0337_),
    .A2(_0332_),
    .A3(_4319_),
    .A4(_4416_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5031_ (.A1(_0469_),
    .A2(_0471_),
    .A3(_0472_),
    .A4(_0473_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5032_ (.A1(_0469_),
    .A2(_0471_),
    .B1(_0472_),
    .B2(_0473_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5033_ (.A1(_0333_),
    .A2(_0373_),
    .A3(_4320_),
    .A4(_0372_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5034_ (.A1(_0371_),
    .A2(_0374_),
    .B(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5035_ (.A1(_0474_),
    .A2(_0475_),
    .A3(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5036_ (.I(_0478_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5037_ (.A1(_0474_),
    .A2(_0475_),
    .B(_0477_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5038_ (.A1(_0463_),
    .A2(_0479_),
    .A3(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5039_ (.A1(_0479_),
    .A2(_0480_),
    .B(_0463_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5040_ (.A1(_0481_),
    .A2(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5041_ (.A1(_0462_),
    .A2(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5042_ (.A1(\as2650.r123[1][3] ),
    .A2(_4304_),
    .B(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5043_ (.A1(_4324_),
    .A2(_0461_),
    .B(_0485_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5044_ (.I(_4325_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5045_ (.A1(\as2650.holding_reg[4] ),
    .A2(_4114_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5046_ (.A1(_4114_),
    .A2(_0425_),
    .B(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5047_ (.A1(_0486_),
    .A2(_0488_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5048_ (.I(\as2650.holding_reg[4] ),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5049_ (.A1(_0419_),
    .A2(_0421_),
    .A3(_0423_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5050_ (.I(_0491_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5051_ (.A1(_0490_),
    .A2(_0492_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5052_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0492_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5053_ (.I(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5054_ (.I(_0407_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5055_ (.A1(_0395_),
    .A2(_0345_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5056_ (.A1(_0384_),
    .A2(_0389_),
    .B1(_0496_),
    .B2(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5057_ (.A1(_0495_),
    .A2(_0498_),
    .B(_0385_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5058_ (.A1(_0495_),
    .A2(_0498_),
    .B(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5059_ (.A1(_0490_),
    .A2(_0426_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5060_ (.A1(_0388_),
    .A2(_0383_),
    .A3(_0392_),
    .B(_0497_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5061_ (.A1(_0501_),
    .A2(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5062_ (.I(_4191_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5063_ (.A1(_0490_),
    .A2(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5064_ (.A1(_4193_),
    .A2(_0427_),
    .B(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5065_ (.A1(_4168_),
    .A2(_0488_),
    .B1(_0506_),
    .B2(_4299_),
    .C(_4165_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5066_ (.A1(_4179_),
    .A2(_0503_),
    .B(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5067_ (.A1(_0410_),
    .A2(_0493_),
    .B1(_0500_),
    .B2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5068_ (.A1(_0489_),
    .A2(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5069_ (.I(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5070_ (.I(_4275_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5071_ (.A1(_0491_),
    .A2(_0448_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5072_ (.A1(_0425_),
    .A2(_0444_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5073_ (.A1(_0512_),
    .A2(_0513_),
    .B1(_0514_),
    .B2(_0455_),
    .C1(_0454_),
    .C2(_0426_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5074_ (.I(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5075_ (.I(_0418_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5076_ (.I(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5077_ (.A1(_4012_),
    .A2(\as2650.r123[1][5] ),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5078_ (.I(\as2650.r123_2[1][5] ),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5079_ (.I(_4019_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5080_ (.A1(_4012_),
    .A2(_0520_),
    .B(_0521_),
    .C(_4002_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5081_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123_2[0][5] ),
    .S(\as2650.psl[4] ),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5082_ (.I(_0523_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5083_ (.I(_0524_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5084_ (.I(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5085_ (.I(_4002_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5086_ (.I(_4019_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5087_ (.A1(_0527_),
    .A2(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5088_ (.A1(_0519_),
    .A2(_0522_),
    .B1(_0526_),
    .B2(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5089_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_4012_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5090_ (.A1(_4213_),
    .A2(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5091_ (.I(\as2650.r0[5] ),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5092_ (.A1(_0533_),
    .A2(_4021_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5093_ (.A1(_0530_),
    .A2(_0532_),
    .A3(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5094_ (.I(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5095_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5096_ (.I(net9),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5097_ (.I(_0538_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5098_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5099_ (.A1(_4042_),
    .A2(_4126_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5100_ (.A1(_0433_),
    .A2(_0345_),
    .B1(_0444_),
    .B2(_0541_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5101_ (.A1(_0492_),
    .A2(_0542_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5102_ (.A1(_4245_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5103_ (.A1(_0540_),
    .A2(_4245_),
    .B(_4227_),
    .C(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5104_ (.A1(_0432_),
    .A2(_0537_),
    .B(_0545_),
    .C(_4204_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5105_ (.A1(_4240_),
    .A2(_0346_),
    .B(_0546_),
    .C(_4198_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5106_ (.A1(_0518_),
    .A2(_4378_),
    .B(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5107_ (.A1(_4369_),
    .A2(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5108_ (.I(_4267_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5109_ (.A1(_0443_),
    .A2(_0425_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5110_ (.A1(_0550_),
    .A2(_0513_),
    .B1(_0514_),
    .B2(_0447_),
    .C(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5111_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5112_ (.A1(_4264_),
    .A2(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5113_ (.A1(_4367_),
    .A2(_0549_),
    .A3(_0554_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5114_ (.A1(_4368_),
    .A2(_0516_),
    .B(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5115_ (.A1(_0292_),
    .A2(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5116_ (.A1(_0293_),
    .A2(_0511_),
    .B(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5117_ (.A1(_0463_),
    .A2(_0478_),
    .A3(_0480_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5118_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123_2[0][4] ),
    .S(\as2650.psl[4] ),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5119_ (.I(_0560_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5120_ (.A1(_4148_),
    .A2(_0561_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5121_ (.I(\as2650.r0[2] ),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5122_ (.I(\as2650.r0[1] ),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5123_ (.A1(_0563_),
    .A2(_0564_),
    .A3(_0368_),
    .A4(_0465_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5124_ (.A1(_4381_),
    .A2(_0368_),
    .B1(_0466_),
    .B2(_4229_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5125_ (.A1(_0565_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5126_ (.A1(_0336_),
    .A2(_4415_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5127_ (.A1(_0417_),
    .A2(_4319_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5128_ (.A1(_0468_),
    .A2(_0568_),
    .A3(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5129_ (.A1(_0562_),
    .A2(_0567_),
    .A3(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5130_ (.I(_0473_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5131_ (.A1(_0572_),
    .A2(_0474_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5132_ (.A1(_0571_),
    .A2(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5133_ (.A1(_0559_),
    .A2(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5134_ (.A1(_0479_),
    .A2(_0574_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5135_ (.A1(_0479_),
    .A2(_0575_),
    .B(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5136_ (.A1(_0462_),
    .A2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5137_ (.A1(\as2650.r123[1][4] ),
    .A2(_4304_),
    .B(_0578_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5138_ (.A1(_4324_),
    .A2(_0558_),
    .B(_0579_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5139_ (.A1(_0323_),
    .A2(_0300_),
    .A3(_0398_),
    .A4(_0424_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5140_ (.A1(_0535_),
    .A2(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5141_ (.A1(_0530_),
    .A2(_0532_),
    .A3(_0534_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5142_ (.A1(_0319_),
    .A2(_0300_),
    .A3(_0398_),
    .A4(_0424_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5143_ (.A1(_0582_),
    .A2(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5144_ (.A1(_4270_),
    .A2(_0535_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5145_ (.A1(_0550_),
    .A2(_0581_),
    .B1(_0584_),
    .B2(_0447_),
    .C(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5146_ (.I(_0586_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5147_ (.I(_0533_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5148_ (.I(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5149_ (.I(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5150_ (.I(_0492_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5151_ (.I(\as2650.r0[6] ),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5152_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5153_ (.A1(_0593_),
    .A2(_4021_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5154_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_4013_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5155_ (.A1(_4214_),
    .A2(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5156_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_4003_),
    .S1(_4013_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5157_ (.A1(_4218_),
    .A2(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5158_ (.A1(_0594_),
    .A2(_0596_),
    .A3(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5159_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5160_ (.I(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5161_ (.I(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5162_ (.I(net1),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5163_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5164_ (.I(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5165_ (.A1(_4077_),
    .A2(_0426_),
    .A3(_0448_),
    .B1(_0583_),
    .B2(_4397_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5166_ (.A1(_0536_),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5167_ (.A1(_0354_),
    .A2(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5168_ (.A1(_0605_),
    .A2(_0354_),
    .B(_0608_),
    .C(_4227_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5169_ (.A1(_0432_),
    .A2(_0602_),
    .B(_0609_),
    .C(_4204_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5170_ (.A1(_4380_),
    .A2(_0591_),
    .B(_0610_),
    .C(_4199_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5171_ (.A1(_0590_),
    .A2(_4378_),
    .B(_4369_),
    .C(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5172_ (.A1(_4370_),
    .A2(_0587_),
    .B(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5173_ (.A1(_4368_),
    .A2(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5174_ (.I(_0582_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5175_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5176_ (.A1(_0322_),
    .A2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5177_ (.A1(_0512_),
    .A2(_0581_),
    .B1(_0584_),
    .B2(_0455_),
    .C(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5178_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5179_ (.A1(_0317_),
    .A2(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5180_ (.A1(_4135_),
    .A2(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5181_ (.I(_0486_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5182_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0616_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5183_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0616_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5184_ (.A1(_0623_),
    .A2(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5185_ (.A1(_0623_),
    .A2(_0624_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5186_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5187_ (.I(_0488_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5188_ (.A1(_0628_),
    .A2(_0493_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5189_ (.A1(_0495_),
    .A2(_0498_),
    .B(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5190_ (.A1(_0627_),
    .A2(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5191_ (.A1(_0385_),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5192_ (.A1(_0495_),
    .A2(_0502_),
    .B(_0493_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5193_ (.A1(_0627_),
    .A2(_0633_),
    .B(_4179_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5194_ (.A1(_0627_),
    .A2(_0633_),
    .B(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5195_ (.I(\as2650.holding_reg[5] ),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5196_ (.A1(_0636_),
    .A2(_4295_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5197_ (.A1(_0396_),
    .A2(_0536_),
    .B(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5198_ (.I(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5199_ (.I(_4193_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5200_ (.I(_0504_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5201_ (.A1(_0636_),
    .A2(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5202_ (.A1(_0640_),
    .A2(_0537_),
    .B(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5203_ (.A1(_0312_),
    .A2(_0639_),
    .B1(_0643_),
    .B2(_0403_),
    .C(_0299_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5204_ (.A1(_0632_),
    .A2(_0635_),
    .A3(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5205_ (.I(_0616_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(_0636_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5207_ (.A1(_0299_),
    .A2(_0647_),
    .B(_0622_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5208_ (.A1(_0622_),
    .A2(_0625_),
    .B1(_0645_),
    .B2(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5209_ (.I(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5210_ (.A1(_0614_),
    .A2(_0621_),
    .B1(_0650_),
    .B2(_4281_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5211_ (.A1(_0571_),
    .A2(_0573_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5212_ (.A1(_0559_),
    .A2(_0574_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5213_ (.A1(_0576_),
    .A2(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5214_ (.A1(_0562_),
    .A2(_0567_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5215_ (.A1(_0655_),
    .A2(_0570_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5216_ (.A1(_0469_),
    .A2(_0568_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5217_ (.A1(_0469_),
    .A2(_0568_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5218_ (.A1(_0657_),
    .A2(_0569_),
    .B(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5219_ (.A1(_0416_),
    .A2(_4414_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5220_ (.A1(_0565_),
    .A2(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5221_ (.A1(_0533_),
    .A2(_4318_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5222_ (.A1(_0661_),
    .A2(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5223_ (.A1(_0562_),
    .A2(_0565_),
    .A3(_0566_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5224_ (.I(\as2650.r0[0] ),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5225_ (.A1(_0564_),
    .A2(_0561_),
    .B1(_0525_),
    .B2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5226_ (.A1(_0564_),
    .A2(_0665_),
    .A3(_0561_),
    .A4(_0525_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5227_ (.A1(_0666_),
    .A2(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5228_ (.A1(_0335_),
    .A2(_0563_),
    .A3(_0367_),
    .A4(_0465_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5229_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5230_ (.A1(_0336_),
    .A2(_0368_),
    .B1(_0466_),
    .B2(_4381_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5231_ (.A1(_0670_),
    .A2(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5232_ (.A1(_0664_),
    .A2(_0668_),
    .A3(_0672_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5233_ (.A1(_0663_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5234_ (.A1(_0656_),
    .A2(_0659_),
    .A3(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5235_ (.A1(_0652_),
    .A2(_0654_),
    .A3(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5236_ (.I(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5237_ (.A1(\as2650.r123[1][5] ),
    .A2(_4413_),
    .B1(_0677_),
    .B2(_4316_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5238_ (.A1(_4138_),
    .A2(_0651_),
    .B(_0678_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5239_ (.A1(_0594_),
    .A2(_0596_),
    .A3(_0598_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5240_ (.I(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5241_ (.I(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5242_ (.A1(\as2650.holding_reg[6] ),
    .A2(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5243_ (.A1(\as2650.holding_reg[6] ),
    .A2(_0599_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5244_ (.A1(_0626_),
    .A2(_0630_),
    .B1(_0638_),
    .B2(_0647_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5245_ (.A1(_0683_),
    .A2(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5246_ (.A1(_0494_),
    .A2(_0502_),
    .B(_0623_),
    .C(_0493_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5247_ (.A1(_0624_),
    .A2(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5248_ (.A1(_0682_),
    .A2(_0687_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5249_ (.I(\as2650.holding_reg[6] ),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5250_ (.A1(_0689_),
    .A2(_0396_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5251_ (.A1(_0396_),
    .A2(_0600_),
    .B(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5252_ (.I(_0691_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5253_ (.A1(_0397_),
    .A2(_0601_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5254_ (.A1(_0689_),
    .A2(_0397_),
    .B(_0403_),
    .C(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5255_ (.A1(_0410_),
    .A2(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5256_ (.A1(_4343_),
    .A2(_0688_),
    .B1(_0692_),
    .B2(_0312_),
    .C(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5257_ (.A1(_4172_),
    .A2(_0685_),
    .B(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(_0689_),
    .A2(_0680_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5259_ (.A1(_0299_),
    .A2(_0698_),
    .B(_0486_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5260_ (.A1(_0622_),
    .A2(_0682_),
    .B1(_0697_),
    .B2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5261_ (.I(_0700_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5262_ (.A1(_4281_),
    .A2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5263_ (.A1(_0615_),
    .A2(_0580_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5264_ (.A1(_0599_),
    .A2(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5265_ (.A1(_0582_),
    .A2(_0583_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5266_ (.A1(_0679_),
    .A2(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5267_ (.A1(_0328_),
    .A2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5268_ (.A1(_0443_),
    .A2(_0600_),
    .B1(_0704_),
    .B2(_0550_),
    .C(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5269_ (.I(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5270_ (.I(_0593_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5271_ (.I(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5272_ (.I(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5273_ (.I(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5274_ (.I(_0537_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5275_ (.A1(_4211_),
    .A2(_4216_),
    .A3(_4220_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5276_ (.I(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5277_ (.I(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5278_ (.A1(_4397_),
    .A2(_0615_),
    .A3(_0583_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5279_ (.A1(_4394_),
    .A2(_0615_),
    .A3(_0580_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5280_ (.A1(_0718_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5281_ (.A1(_0601_),
    .A2(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5282_ (.A1(_4247_),
    .A2(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5283_ (.I(net2),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5284_ (.I(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5285_ (.I(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5286_ (.I(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5287_ (.A1(_0726_),
    .A2(_4247_),
    .B(_4252_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5288_ (.A1(_0432_),
    .A2(_0717_),
    .B1(_0722_),
    .B2(_0727_),
    .C(_4204_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5289_ (.A1(_4380_),
    .A2(_0714_),
    .B(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5290_ (.A1(_4378_),
    .A2(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5291_ (.A1(_0713_),
    .A2(_4201_),
    .B(_4258_),
    .C(_0730_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5292_ (.A1(_4370_),
    .A2(_0709_),
    .B(_0731_),
    .C(_0317_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5293_ (.A1(_0318_),
    .A2(_0706_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5294_ (.A1(_0454_),
    .A2(_0600_),
    .B1(_0704_),
    .B2(_0512_),
    .C(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5295_ (.I(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(_4280_),
    .A2(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5297_ (.A1(_0293_),
    .A2(_0732_),
    .A3(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5298_ (.A1(_0702_),
    .A2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(_0652_),
    .A2(_0675_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5300_ (.A1(_0652_),
    .A2(_0675_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5301_ (.A1(_0654_),
    .A2(_0739_),
    .B(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5302_ (.A1(_0656_),
    .A2(_0674_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5303_ (.A1(_0656_),
    .A2(_0674_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5304_ (.A1(_0659_),
    .A2(_0742_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5305_ (.A1(_0418_),
    .A2(_0372_),
    .A3(_0565_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5306_ (.A1(_0661_),
    .A2(_0662_),
    .B(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5307_ (.A1(_0666_),
    .A2(_0667_),
    .A3(_0670_),
    .A4(_0671_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5308_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_0670_),
    .B2(_0671_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5309_ (.A1(_0664_),
    .A2(_0747_),
    .A3(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5310_ (.A1(_0663_),
    .A2(_0673_),
    .B(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5311_ (.I(\as2650.r0[5] ),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5312_ (.A1(_0751_),
    .A2(_4415_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5313_ (.A1(_0669_),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5314_ (.A1(_0593_),
    .A2(_4318_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5315_ (.A1(_0753_),
    .A2(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5316_ (.A1(_0336_),
    .A2(_0467_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5317_ (.A1(_0417_),
    .A2(_0369_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5318_ (.A1(_0335_),
    .A2(_0367_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(\as2650.r0[4] ),
    .A2(_0464_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5320_ (.A1(_0758_),
    .A2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5321_ (.A1(_0756_),
    .A2(_0757_),
    .B(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5322_ (.A1(\as2650.r0[1] ),
    .A2(_0523_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5323_ (.A1(\as2650.r0[2] ),
    .A2(_0560_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5324_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .S(\as2650.psl[4] ),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5325_ (.I(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5326_ (.A1(\as2650.r0[0] ),
    .A2(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5327_ (.A1(_0762_),
    .A2(_0763_),
    .A3(_0766_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5328_ (.A1(_0667_),
    .A2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5329_ (.A1(_0747_),
    .A2(_0761_),
    .A3(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5330_ (.A1(_0750_),
    .A2(_0755_),
    .A3(_0769_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5331_ (.A1(_0746_),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5332_ (.A1(_0744_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5333_ (.A1(_0741_),
    .A2(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5334_ (.I(_0773_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5335_ (.A1(\as2650.r123[1][6] ),
    .A2(_4413_),
    .B1(_0774_),
    .B2(_4316_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5336_ (.A1(_4138_),
    .A2(_0738_),
    .B(_0775_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5337_ (.A1(_0680_),
    .A2(_0703_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5338_ (.A1(_0715_),
    .A2(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5339_ (.A1(_0599_),
    .A2(_0705_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5340_ (.A1(_0715_),
    .A2(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5341_ (.A1(_4222_),
    .A2(_0443_),
    .B1(_0777_),
    .B2(_0550_),
    .C1(_0779_),
    .C2(_0447_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5342_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5343_ (.A1(_4206_),
    .A2(_4379_),
    .B(_4174_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5344_ (.I(net3),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5345_ (.I(_0783_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5346_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5347_ (.I0(_0718_),
    .I1(_0719_),
    .S(_0679_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5348_ (.A1(_4221_),
    .A2(_0786_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5349_ (.A1(_4246_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5350_ (.A1(_0785_),
    .A2(_4246_),
    .B(_4228_),
    .C(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5351_ (.A1(_4228_),
    .A2(_0782_),
    .B(_0789_),
    .C(_4205_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5352_ (.A1(_4205_),
    .A2(_0681_),
    .B(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5353_ (.I(_4210_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5354_ (.A1(_0792_),
    .A2(_4200_),
    .B(_4258_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5355_ (.A1(_4200_),
    .A2(_0791_),
    .B(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5356_ (.A1(_4264_),
    .A2(_0781_),
    .B(_0794_),
    .C(_4280_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5357_ (.A1(_4222_),
    .A2(_0454_),
    .B1(_0777_),
    .B2(_0512_),
    .C1(_0779_),
    .C2(_0455_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5358_ (.I(_0796_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5359_ (.A1(_4368_),
    .A2(_0797_),
    .B(_0293_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5360_ (.I(\as2650.holding_reg[7] ),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5361_ (.A1(_0799_),
    .A2(_4222_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5362_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0716_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5363_ (.A1(_0800_),
    .A2(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5364_ (.I(_0802_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5365_ (.A1(_0622_),
    .A2(_0803_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5366_ (.A1(_0698_),
    .A2(_0691_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5367_ (.A1(_0682_),
    .A2(_0684_),
    .B(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5368_ (.A1(_0802_),
    .A2(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5369_ (.A1(_0624_),
    .A2(_0683_),
    .A3(_0686_),
    .B(_0698_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5370_ (.A1(_0802_),
    .A2(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5371_ (.A1(_0799_),
    .A2(_0641_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5372_ (.A1(_0641_),
    .A2(_0716_),
    .B(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5373_ (.A1(_4179_),
    .A2(_0809_),
    .B1(_0811_),
    .B2(_4171_),
    .C(_4348_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5374_ (.A1(_0385_),
    .A2(_0807_),
    .B(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5375_ (.A1(_0405_),
    .A2(_0800_),
    .B(_4164_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _5376_ (.A1(_0410_),
    .A2(_0801_),
    .B1(_0813_),
    .B2(_0814_),
    .C(_4147_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5377_ (.A1(_4139_),
    .A2(_0804_),
    .A3(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5378_ (.A1(_0795_),
    .A2(_0798_),
    .B(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5379_ (.I(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5380_ (.A1(_0744_),
    .A2(_0771_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5381_ (.A1(_0741_),
    .A2(_0772_),
    .B(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5382_ (.A1(_0747_),
    .A2(_0761_),
    .A3(_0768_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5383_ (.A1(_0755_),
    .A2(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5384_ (.A1(_0755_),
    .A2(_0821_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5385_ (.A1(_0750_),
    .A2(_0822_),
    .A3(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5386_ (.A1(_0746_),
    .A2(_0770_),
    .B(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5387_ (.A1(_0588_),
    .A2(_4417_),
    .A3(_0670_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5388_ (.A1(_0710_),
    .A2(_4321_),
    .A3(_0753_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5389_ (.A1(_0826_),
    .A2(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5390_ (.A1(_0761_),
    .A2(_0768_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5391_ (.A1(_0668_),
    .A2(_0672_),
    .A3(_0829_),
    .B1(_0821_),
    .B2(_0755_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5392_ (.A1(\as2650.r0[6] ),
    .A2(_4414_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5393_ (.A1(_0760_),
    .A2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5394_ (.A1(\as2650.r0[7] ),
    .A2(_4318_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5395_ (.A1(_0832_),
    .A2(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5396_ (.A1(_0562_),
    .A2(_0762_),
    .A3(_0767_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5397_ (.A1(_0761_),
    .A2(_0768_),
    .B(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5398_ (.I(_0759_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5399_ (.A1(\as2650.r0[5] ),
    .A2(_0367_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5400_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_4009_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5401_ (.A1(_4148_),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5402_ (.A1(_0837_),
    .A2(_0838_),
    .A3(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5403_ (.I(_0524_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5404_ (.A1(_0665_),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5405_ (.A1(\as2650.r0[1] ),
    .A2(_0764_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5406_ (.I(_0765_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5407_ (.A1(_0564_),
    .A2(_0525_),
    .B1(_0845_),
    .B2(_0665_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5408_ (.A1(_0843_),
    .A2(_0844_),
    .B1(_0846_),
    .B2(_0763_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5409_ (.A1(\as2650.r0[3] ),
    .A2(_0560_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5410_ (.A1(_0563_),
    .A2(_0524_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5411_ (.A1(_0844_),
    .A2(_0848_),
    .A3(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5412_ (.A1(_0847_),
    .A2(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5413_ (.A1(_0841_),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5414_ (.A1(_0834_),
    .A2(_0836_),
    .A3(_0852_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5415_ (.A1(_0830_),
    .A2(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5416_ (.A1(_0828_),
    .A2(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5417_ (.A1(_0825_),
    .A2(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5418_ (.A1(_0820_),
    .A2(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5419_ (.A1(_4302_),
    .A2(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5420_ (.A1(\as2650.r123[1][7] ),
    .A2(_4304_),
    .B(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5421_ (.A1(_4138_),
    .A2(_0818_),
    .B(_0859_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5422_ (.I(_0528_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5423_ (.I(_4110_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5424_ (.A1(_4111_),
    .A2(_4086_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5425_ (.A1(_4111_),
    .A2(_0353_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5426_ (.A1(_4361_),
    .A2(_4096_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5427_ (.A1(_4093_),
    .A2(_4091_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5428_ (.A1(_4111_),
    .A2(_0864_),
    .A3(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5429_ (.A1(_0862_),
    .A2(_0863_),
    .A3(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5430_ (.A1(_0861_),
    .A2(_0867_),
    .B(_4134_),
    .C(_4117_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5431_ (.A1(_0860_),
    .A2(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5432_ (.I(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5433_ (.I(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5434_ (.A1(_4004_),
    .A2(_0521_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5435_ (.A1(_0504_),
    .A2(_4299_),
    .A3(_4300_),
    .A4(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5436_ (.A1(_4067_),
    .A2(_4144_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5437_ (.A1(_4163_),
    .A2(_4296_),
    .A3(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5438_ (.A1(_0873_),
    .A2(_0875_),
    .B(_4291_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5439_ (.A1(_4017_),
    .A2(_0876_),
    .B(_0870_),
    .C(_4285_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5440_ (.I(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5441_ (.I(_0875_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5442_ (.I(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5443_ (.I(_0880_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5444_ (.I(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5445_ (.I(_4109_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5446_ (.A1(_4140_),
    .A2(_0874_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5447_ (.A1(_4311_),
    .A2(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5448_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5449_ (.I(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5450_ (.A1(_0883_),
    .A2(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5451_ (.A1(_4290_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5452_ (.I(\as2650.psu[0] ),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5453_ (.A1(_0890_),
    .A2(\as2650.psu[1] ),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5454_ (.I(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5455_ (.I(_0892_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5456_ (.I(\as2650.psu[0] ),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5457_ (.I(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5458_ (.I(\as2650.psu[1] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5460_ (.A1(_0895_),
    .A2(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5461_ (.I(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5462_ (.I(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5463_ (.A1(\as2650.stack[3][8] ),
    .A2(_0893_),
    .B1(_0900_),
    .B2(\as2650.stack[2][8] ),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5464_ (.I(\as2650.psu[1] ),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5465_ (.A1(_0895_),
    .A2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5466_ (.I(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5467_ (.I(_0890_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5468_ (.A1(_0905_),
    .A2(_0897_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5469_ (.I(_0906_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5470_ (.I(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5471_ (.A1(\as2650.psu[2] ),
    .A2(_0891_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5472_ (.I(\as2650.psu[2] ),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5473_ (.A1(_0894_),
    .A2(_0896_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5474_ (.A1(_0910_),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5475_ (.A1(_0909_),
    .A2(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5476_ (.I(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5477_ (.I(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5478_ (.I(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5479_ (.A1(\as2650.stack[0][8] ),
    .A2(_0904_),
    .B1(_0908_),
    .B2(\as2650.stack[1][8] ),
    .C(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5480_ (.I(_0907_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5481_ (.A1(\as2650.stack[4][8] ),
    .A2(_0904_),
    .B1(_0918_),
    .B2(\as2650.stack[5][8] ),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5482_ (.I(_0898_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5483_ (.A1(_0909_),
    .A2(_0912_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5484_ (.I(_0921_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5485_ (.I(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5486_ (.A1(\as2650.stack[7][8] ),
    .A2(_0893_),
    .B1(_0920_),
    .B2(\as2650.stack[6][8] ),
    .C(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5487_ (.A1(_0901_),
    .A2(_0917_),
    .B1(_0919_),
    .B2(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5488_ (.A1(_4129_),
    .A2(_4312_),
    .A3(_0529_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5489_ (.A1(_4313_),
    .A2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5490_ (.A1(_0879_),
    .A2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5491_ (.A1(_4309_),
    .A2(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5492_ (.I(_0929_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5493_ (.A1(_4306_),
    .A2(_0882_),
    .B1(_0889_),
    .B2(_0925_),
    .C(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5494_ (.A1(_4283_),
    .A2(_0871_),
    .B(_0878_),
    .C(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5495_ (.I(\as2650.r123[0][0] ),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5496_ (.I(_0926_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5497_ (.I(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5498_ (.I(_0886_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5499_ (.I(_4108_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5500_ (.I(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5501_ (.A1(_0935_),
    .A2(_0936_),
    .B(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5502_ (.I(net10),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5503_ (.A1(_4290_),
    .A2(_0939_),
    .B(_0869_),
    .C(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5504_ (.I(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5505_ (.A1(_0933_),
    .A2(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5506_ (.A1(_0932_),
    .A2(_0943_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5507_ (.I(_0944_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5508_ (.I(_0860_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5509_ (.I(_0941_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5510_ (.I(_0881_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5511_ (.I(_0909_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5512_ (.I(_0912_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5513_ (.I(_0949_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5514_ (.A1(\as2650.stack[3][9] ),
    .A2(_0948_),
    .B(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5515_ (.I(_0898_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5516_ (.I(_0903_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5517_ (.A1(\as2650.stack[0][9] ),
    .A2(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5518_ (.A1(\as2650.stack[2][9] ),
    .A2(_0952_),
    .B1(_0908_),
    .B2(\as2650.stack[1][9] ),
    .C(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5519_ (.A1(\as2650.stack[4][9] ),
    .A2(_0904_),
    .B1(_0918_),
    .B2(\as2650.stack[5][9] ),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5520_ (.I(_0923_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5521_ (.A1(\as2650.stack[7][9] ),
    .A2(_0893_),
    .B1(_0952_),
    .B2(\as2650.stack[6][9] ),
    .C(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5522_ (.A1(_0951_),
    .A2(_0955_),
    .B1(_0956_),
    .B2(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5523_ (.A1(_4377_),
    .A2(_0947_),
    .B1(_0889_),
    .B2(_0959_),
    .C(_0929_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5524_ (.A1(_0946_),
    .A2(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5525_ (.A1(\as2650.r123[0][1] ),
    .A2(_0942_),
    .B(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5526_ (.A1(_0945_),
    .A2(_4136_),
    .A3(_4412_),
    .B(_0962_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5527_ (.I(_0877_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5528_ (.A1(\as2650.r123[0][2] ),
    .A2(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5529_ (.A1(_4308_),
    .A2(_0880_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5530_ (.A1(_4017_),
    .A2(_0965_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5531_ (.I(_0909_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5532_ (.A1(\as2650.stack[3][10] ),
    .A2(_0967_),
    .B(_0950_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5533_ (.I(_0899_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5534_ (.A1(\as2650.stack[2][10] ),
    .A2(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5535_ (.I(_0953_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5536_ (.I(_0906_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5537_ (.I(_0972_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5538_ (.A1(\as2650.stack[0][10] ),
    .A2(_0971_),
    .B1(_0973_),
    .B2(\as2650.stack[1][10] ),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5539_ (.A1(_0968_),
    .A2(_0970_),
    .A3(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5540_ (.A1(\as2650.stack[4][10] ),
    .A2(_0971_),
    .B1(_0973_),
    .B2(\as2650.stack[5][10] ),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5541_ (.I(_0892_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5542_ (.A1(\as2650.stack[7][10] ),
    .A2(_0977_),
    .B1(_0969_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5543_ (.A1(_0916_),
    .A2(_0976_),
    .A3(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5544_ (.A1(_0975_),
    .A2(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5545_ (.I(_0334_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5546_ (.A1(_0981_),
    .A2(_0947_),
    .B(_0929_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5547_ (.A1(_0966_),
    .A2(_0980_),
    .B(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5548_ (.A1(_0366_),
    .A2(_0870_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5549_ (.A1(_0946_),
    .A2(_0983_),
    .A3(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5550_ (.A1(_0964_),
    .A2(_0985_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5551_ (.A1(\as2650.r123[0][3] ),
    .A2(_0878_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5552_ (.A1(\as2650.stack[3][11] ),
    .A2(_0948_),
    .B(_0950_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5553_ (.I(_0903_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5554_ (.A1(\as2650.stack[1][11] ),
    .A2(_0972_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5555_ (.A1(\as2650.stack[2][11] ),
    .A2(_0920_),
    .B1(_0988_),
    .B2(\as2650.stack[0][11] ),
    .C(_0989_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5556_ (.A1(\as2650.stack[7][11] ),
    .A2(_0891_),
    .B1(_0903_),
    .B2(\as2650.stack[4][11] ),
    .C1(\as2650.stack[5][11] ),
    .C2(_0907_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5557_ (.A1(_0915_),
    .A2(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5558_ (.A1(\as2650.stack[6][11] ),
    .A2(_0952_),
    .B(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5559_ (.A1(_0987_),
    .A2(_0990_),
    .B(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5560_ (.A1(_0415_),
    .A2(_0882_),
    .B1(_0889_),
    .B2(_0994_),
    .C(_0930_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5561_ (.A1(_0461_),
    .A2(_0871_),
    .B(_0963_),
    .C(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5562_ (.A1(_0986_),
    .A2(_0996_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5563_ (.I(_0997_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5564_ (.I(\as2650.r123[0][4] ),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5565_ (.A1(_0998_),
    .A2(_0942_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5566_ (.I(_0517_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5567_ (.A1(\as2650.stack[3][12] ),
    .A2(_0948_),
    .B(_0949_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5568_ (.A1(\as2650.stack[2][12] ),
    .A2(_0920_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5569_ (.A1(\as2650.stack[0][12] ),
    .A2(_0953_),
    .B1(_0972_),
    .B2(\as2650.stack[1][12] ),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5570_ (.A1(_1001_),
    .A2(_1002_),
    .A3(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5571_ (.A1(\as2650.stack[4][12] ),
    .A2(_0988_),
    .B1(_0972_),
    .B2(\as2650.stack[5][12] ),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5572_ (.A1(\as2650.stack[7][12] ),
    .A2(_0892_),
    .B1(_0899_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5573_ (.A1(_0916_),
    .A2(_1005_),
    .A3(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5574_ (.A1(_1004_),
    .A2(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5575_ (.A1(_0966_),
    .A2(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5576_ (.A1(_1000_),
    .A2(_0966_),
    .B(_0930_),
    .C(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5577_ (.A1(_0558_),
    .A2(_0871_),
    .B(_0963_),
    .C(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5578_ (.A1(_0999_),
    .A2(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5579_ (.I(_1012_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5580_ (.I(\as2650.r123[0][5] ),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5581_ (.A1(\as2650.stack[3][13] ),
    .A2(_0948_),
    .B(_0950_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5582_ (.A1(\as2650.stack[2][13] ),
    .A2(_0969_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5583_ (.A1(\as2650.stack[0][13] ),
    .A2(_0904_),
    .B1(_0918_),
    .B2(\as2650.stack[1][13] ),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5584_ (.A1(_1014_),
    .A2(_1015_),
    .A3(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5585_ (.A1(\as2650.stack[4][13] ),
    .A2(_0971_),
    .B1(_0918_),
    .B2(\as2650.stack[5][13] ),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5586_ (.A1(\as2650.stack[7][13] ),
    .A2(_0977_),
    .B1(_0900_),
    .B2(\as2650.stack[6][13] ),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5587_ (.A1(_0916_),
    .A2(_1018_),
    .A3(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5588_ (.A1(_1017_),
    .A2(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5589_ (.I(_0589_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5590_ (.A1(_1022_),
    .A2(_0947_),
    .B(_0929_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5591_ (.A1(_0966_),
    .A2(_1021_),
    .B(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5592_ (.A1(_0651_),
    .A2(_0870_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5593_ (.A1(_0946_),
    .A2(_1024_),
    .A3(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5594_ (.A1(_1013_),
    .A2(_0942_),
    .B(_1026_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5595_ (.A1(\as2650.r123[0][6] ),
    .A2(_0878_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5596_ (.I(_0711_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5597_ (.A1(\as2650.stack[6][14] ),
    .A2(_0952_),
    .B1(_0988_),
    .B2(\as2650.stack[4][14] ),
    .C1(\as2650.stack[5][14] ),
    .C2(_0908_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5598_ (.A1(\as2650.stack[7][14] ),
    .A2(_0977_),
    .B(_0957_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5599_ (.A1(\as2650.stack[0][14] ),
    .A2(_0953_),
    .B1(_0907_),
    .B2(\as2650.stack[1][14] ),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5600_ (.I(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5601_ (.A1(\as2650.stack[3][14] ),
    .A2(_0893_),
    .B1(_0900_),
    .B2(\as2650.stack[2][14] ),
    .C(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5602_ (.A1(_1029_),
    .A2(_1030_),
    .B1(_1033_),
    .B2(_0957_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5603_ (.A1(_1028_),
    .A2(_0882_),
    .B1(_0889_),
    .B2(_1034_),
    .C(_0930_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5604_ (.A1(_0738_),
    .A2(_0871_),
    .B(_0878_),
    .C(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5605_ (.A1(_1027_),
    .A2(_1036_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5606_ (.I(_1037_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5607_ (.A1(\as2650.r123[0][7] ),
    .A2(_0963_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5608_ (.I(_0792_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5609_ (.I(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5610_ (.A1(_1040_),
    .A2(_4309_),
    .A3(_0882_),
    .A4(_0928_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5611_ (.A1(_0817_),
    .A2(_0869_),
    .B(_0946_),
    .C(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5612_ (.A1(_1038_),
    .A2(_1042_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5613_ (.I(\as2650.psu[2] ),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5614_ (.I(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5615_ (.A1(_0890_),
    .A2(_0902_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5616_ (.I(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5617_ (.I(_1046_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5618_ (.I(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5619_ (.A1(_4141_),
    .A2(_0504_),
    .A3(_0872_),
    .A4(_0874_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5620_ (.A1(_4038_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5621_ (.A1(_4288_),
    .A2(_1050_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5622_ (.I(_0351_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5623_ (.I(\as2650.cycle[2] ),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5624_ (.I(_1053_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5625_ (.A1(_4029_),
    .A2(_1054_),
    .A3(_4119_),
    .A4(_4033_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5626_ (.A1(_4102_),
    .A2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5627_ (.I(_4118_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5628_ (.I(_4120_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5629_ (.A1(_4050_),
    .A2(\as2650.cycle[4] ),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5630_ (.A1(_4046_),
    .A2(_4051_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5631_ (.A1(_1059_),
    .A2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5632_ (.A1(_1058_),
    .A2(_4121_),
    .A3(_4119_),
    .A4(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5633_ (.A1(_1057_),
    .A2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5634_ (.A1(_1056_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5635_ (.A1(\as2650.addr_buff[7] ),
    .A2(_4124_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5636_ (.A1(_1064_),
    .A2(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5637_ (.A1(_1052_),
    .A2(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5638_ (.A1(_4163_),
    .A2(_4089_),
    .A3(_4074_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5639_ (.I(_4080_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5640_ (.A1(_4170_),
    .A2(_4044_),
    .A3(_4214_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5641_ (.A1(_1069_),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5642_ (.I(_4124_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5643_ (.I(_4063_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5644_ (.I(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5645_ (.A1(\as2650.ins_reg[3] ),
    .A2(_4067_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5646_ (.A1(_4003_),
    .A2(_0528_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5647_ (.A1(_4297_),
    .A2(_1075_),
    .A3(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5648_ (.I(_1077_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5649_ (.A1(_1074_),
    .A2(_1078_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5650_ (.A1(_4142_),
    .A2(_1072_),
    .A3(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5651_ (.A1(_1067_),
    .A2(_1068_),
    .A3(_1071_),
    .B(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5652_ (.A1(_4110_),
    .A2(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5653_ (.A1(_1051_),
    .A2(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5654_ (.I(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5655_ (.A1(_1044_),
    .A2(_1048_),
    .A3(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5656_ (.I(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5657_ (.I(_1086_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5658_ (.I(\as2650.pc[8] ),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5659_ (.I(_1051_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5660_ (.I(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5661_ (.I(_4083_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5662_ (.A1(_4129_),
    .A2(_0529_),
    .A3(_0884_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5663_ (.A1(_1091_),
    .A2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5664_ (.I(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5665_ (.A1(_4015_),
    .A2(_4288_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5666_ (.I(_1095_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5667_ (.A1(_1094_),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5668_ (.I(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5669_ (.I(_4289_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5670_ (.I(_1094_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5671_ (.A1(_0933_),
    .A2(_1099_),
    .A3(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5672_ (.A1(_1088_),
    .A2(_1090_),
    .B1(_1098_),
    .B2(\as2650.r123_2[0][0] ),
    .C(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5673_ (.I(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5674_ (.I(_1086_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5675_ (.A1(\as2650.stack[3][8] ),
    .A2(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5676_ (.A1(_1087_),
    .A2(_1103_),
    .B(_1105_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5677_ (.I(\as2650.pc[9] ),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5678_ (.I(\as2650.r123[0][1] ),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5679_ (.A1(_1107_),
    .A2(_1099_),
    .A3(_1100_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5680_ (.A1(_1106_),
    .A2(_1090_),
    .B1(_1098_),
    .B2(\as2650.r123_2[0][1] ),
    .C(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5681_ (.I(_1109_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5682_ (.I(_1085_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5683_ (.A1(\as2650.stack[3][9] ),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5684_ (.A1(_1087_),
    .A2(_1110_),
    .B(_1112_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5685_ (.A1(_1099_),
    .A2(_1100_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5686_ (.I(\as2650.pc[10] ),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5687_ (.A1(_1114_),
    .A2(_1089_),
    .B1(_1097_),
    .B2(\as2650.r123_2[0][2] ),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5688_ (.I(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5689_ (.A1(\as2650.r123[0][2] ),
    .A2(_1113_),
    .B(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5690_ (.I(_1117_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5691_ (.A1(\as2650.stack[3][10] ),
    .A2(_1111_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5692_ (.A1(_1087_),
    .A2(_1118_),
    .B(_1119_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5693_ (.I(\as2650.pc[11] ),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5695_ (.I(_1121_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5696_ (.A1(_1122_),
    .A2(_1089_),
    .B1(_1097_),
    .B2(\as2650.r123_2[0][3] ),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5697_ (.I(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5698_ (.A1(\as2650.r123[0][3] ),
    .A2(_1113_),
    .B(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5699_ (.I(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5700_ (.A1(\as2650.stack[3][11] ),
    .A2(_1111_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5701_ (.A1(_1087_),
    .A2(_1126_),
    .B(_1127_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5702_ (.I(\as2650.pc[12] ),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5703_ (.I(_1128_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5704_ (.I(_1129_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5705_ (.A1(_0998_),
    .A2(_1099_),
    .A3(_1100_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5706_ (.A1(_1130_),
    .A2(_1090_),
    .B1(_1098_),
    .B2(\as2650.r123_2[0][4] ),
    .C(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5707_ (.I(_1132_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5708_ (.A1(\as2650.stack[3][12] ),
    .A2(_1111_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5709_ (.A1(_1104_),
    .A2(_1133_),
    .B(_1134_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5710_ (.I(\as2650.pc[13] ),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5711_ (.A1(_1013_),
    .A2(_4290_),
    .A3(_1094_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5712_ (.A1(_1135_),
    .A2(_1090_),
    .B1(_1098_),
    .B2(\as2650.r123_2[0][5] ),
    .C(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5713_ (.I(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5714_ (.A1(\as2650.stack[3][13] ),
    .A2(_1086_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5715_ (.A1(_1104_),
    .A2(_1138_),
    .B(_1139_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5716_ (.A1(\as2650.pc[14] ),
    .A2(_1089_),
    .B1(_1097_),
    .B2(\as2650.r123_2[0][6] ),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5717_ (.I(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5718_ (.A1(\as2650.r123[0][6] ),
    .A2(_1113_),
    .B(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5719_ (.I(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5720_ (.A1(\as2650.stack[3][14] ),
    .A2(_1086_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5721_ (.A1(_1104_),
    .A2(_1143_),
    .B(_1144_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5722_ (.I(_1083_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5723_ (.I(_1043_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5724_ (.A1(_1146_),
    .A2(_0988_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5725_ (.A1(_1145_),
    .A2(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5726_ (.I(_1148_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5727_ (.I(_1149_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5728_ (.I(_1149_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5729_ (.A1(\as2650.stack[5][8] ),
    .A2(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5730_ (.A1(_1103_),
    .A2(_1150_),
    .B(_1152_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5731_ (.I(_1148_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5732_ (.A1(\as2650.stack[5][9] ),
    .A2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5733_ (.A1(_1110_),
    .A2(_1150_),
    .B(_1154_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5734_ (.A1(\as2650.stack[5][10] ),
    .A2(_1153_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5735_ (.A1(_1118_),
    .A2(_1150_),
    .B(_1155_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5736_ (.A1(\as2650.stack[5][11] ),
    .A2(_1153_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5737_ (.A1(_1126_),
    .A2(_1150_),
    .B(_1156_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5738_ (.A1(\as2650.stack[5][12] ),
    .A2(_1153_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5739_ (.A1(_1133_),
    .A2(_1151_),
    .B(_1157_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5740_ (.A1(\as2650.stack[5][13] ),
    .A2(_1149_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5741_ (.A1(_1138_),
    .A2(_1151_),
    .B(_1158_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5742_ (.A1(\as2650.stack[5][14] ),
    .A2(_1149_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5743_ (.A1(_1143_),
    .A2(_1151_),
    .B(_1159_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5744_ (.A1(_1146_),
    .A2(_0908_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5745_ (.A1(_1145_),
    .A2(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5746_ (.I(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5747_ (.I(_1162_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5748_ (.I(_1162_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5749_ (.A1(\as2650.stack[6][8] ),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5750_ (.A1(_1103_),
    .A2(_1163_),
    .B(_1165_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5751_ (.I(_1161_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5752_ (.A1(\as2650.stack[6][9] ),
    .A2(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5753_ (.A1(_1110_),
    .A2(_1163_),
    .B(_1167_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5754_ (.A1(\as2650.stack[6][10] ),
    .A2(_1166_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5755_ (.A1(_1118_),
    .A2(_1163_),
    .B(_1168_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5756_ (.A1(\as2650.stack[6][11] ),
    .A2(_1166_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5757_ (.A1(_1126_),
    .A2(_1163_),
    .B(_1169_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5758_ (.A1(\as2650.stack[6][12] ),
    .A2(_1166_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5759_ (.A1(_1133_),
    .A2(_1164_),
    .B(_1170_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5760_ (.A1(\as2650.stack[6][13] ),
    .A2(_1162_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5761_ (.A1(_1138_),
    .A2(_1164_),
    .B(_1171_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5762_ (.A1(\as2650.stack[6][14] ),
    .A2(_1162_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5763_ (.A1(_1143_),
    .A2(_1164_),
    .B(_1172_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5764_ (.I(_1043_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5765_ (.I(_1173_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5766_ (.A1(_0895_),
    .A2(\as2650.psu[1] ),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5767_ (.I(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5768_ (.I(_1176_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5769_ (.A1(_1174_),
    .A2(_1177_),
    .A3(_1084_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5770_ (.I(_1178_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5771_ (.I(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5772_ (.I(_1179_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5773_ (.A1(\as2650.stack[2][8] ),
    .A2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5774_ (.A1(_1103_),
    .A2(_1180_),
    .B(_1182_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5775_ (.I(_1178_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5776_ (.A1(\as2650.stack[2][9] ),
    .A2(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5777_ (.A1(_1110_),
    .A2(_1180_),
    .B(_1184_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5778_ (.A1(\as2650.stack[2][10] ),
    .A2(_1183_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5779_ (.A1(_1118_),
    .A2(_1180_),
    .B(_1185_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5780_ (.A1(\as2650.stack[2][11] ),
    .A2(_1183_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5781_ (.A1(_1126_),
    .A2(_1180_),
    .B(_1186_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5782_ (.A1(\as2650.stack[2][12] ),
    .A2(_1183_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5783_ (.A1(_1133_),
    .A2(_1181_),
    .B(_1187_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5784_ (.A1(\as2650.stack[2][13] ),
    .A2(_1179_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5785_ (.A1(_1138_),
    .A2(_1181_),
    .B(_1188_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5786_ (.A1(\as2650.stack[2][14] ),
    .A2(_1179_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5787_ (.A1(_1143_),
    .A2(_1181_),
    .B(_1189_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5788_ (.I(_1102_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5789_ (.A1(_0890_),
    .A2(_0897_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5790_ (.I(_1191_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5791_ (.I(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5792_ (.I(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5793_ (.A1(_1044_),
    .A2(_1194_),
    .A3(_1084_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5794_ (.I(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5795_ (.I(_1196_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5796_ (.I(_1196_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5797_ (.A1(\as2650.stack[1][8] ),
    .A2(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5798_ (.A1(_1190_),
    .A2(_1197_),
    .B(_1199_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5799_ (.I(_1109_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5800_ (.I(_1195_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5801_ (.A1(\as2650.stack[1][9] ),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5802_ (.A1(_1200_),
    .A2(_1197_),
    .B(_1202_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5803_ (.I(_1117_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5804_ (.A1(\as2650.stack[1][10] ),
    .A2(_1201_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5805_ (.A1(_1203_),
    .A2(_1197_),
    .B(_1204_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5806_ (.I(_1125_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5807_ (.A1(\as2650.stack[1][11] ),
    .A2(_1201_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5808_ (.A1(_1205_),
    .A2(_1197_),
    .B(_1206_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5809_ (.I(_1132_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5810_ (.A1(\as2650.stack[1][12] ),
    .A2(_1201_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5811_ (.A1(_1207_),
    .A2(_1198_),
    .B(_1208_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5812_ (.I(_1137_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5813_ (.A1(\as2650.stack[1][13] ),
    .A2(_1196_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5814_ (.A1(_1209_),
    .A2(_1198_),
    .B(_1210_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5815_ (.I(_1142_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5816_ (.A1(\as2650.stack[1][14] ),
    .A2(_1196_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5817_ (.A1(_1211_),
    .A2(_1198_),
    .B(_1212_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5818_ (.I(\as2650.psu[5] ),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5819_ (.I(_4307_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5820_ (.A1(_4314_),
    .A2(_0926_),
    .A3(_0885_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5821_ (.A1(_0860_),
    .A2(_4295_),
    .A3(_4312_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5822_ (.I(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5823_ (.A1(_0860_),
    .A2(_4295_),
    .A3(_0884_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5824_ (.I(_1218_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5825_ (.A1(_4006_),
    .A2(_1217_),
    .B(_1219_),
    .C(_1092_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5826_ (.A1(_1215_),
    .A2(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5827_ (.A1(_1073_),
    .A2(_4099_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5828_ (.I(_1222_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5829_ (.I(_4073_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5830_ (.A1(_1224_),
    .A2(_4128_),
    .A3(_4145_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5831_ (.A1(_1223_),
    .A2(_1225_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5832_ (.A1(_4079_),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5833_ (.A1(_1214_),
    .A2(_1221_),
    .A3(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5834_ (.A1(_1073_),
    .A2(_4087_),
    .A3(_4144_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5835_ (.I(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5836_ (.I(_0405_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5837_ (.I(_4214_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5838_ (.A1(\as2650.psl[6] ),
    .A2(_4004_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5839_ (.A1(\as2650.psl[7] ),
    .A2(_0528_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5840_ (.A1(_1233_),
    .A2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5841_ (.A1(_1232_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5842_ (.A1(_0938_),
    .A2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5843_ (.A1(_1231_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5844_ (.A1(_1230_),
    .A2(_1238_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5845_ (.I(_1074_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5846_ (.I(_4040_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5847_ (.I(_1241_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5848_ (.I(_4027_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5849_ (.A1(_1240_),
    .A2(_1242_),
    .A3(_1243_),
    .A4(_0350_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5850_ (.I(_1244_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5851_ (.A1(_1058_),
    .A2(_1053_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5852_ (.A1(_4032_),
    .A2(_4118_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5853_ (.A1(_1061_),
    .A2(_1246_),
    .A3(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5854_ (.I(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5855_ (.A1(_1232_),
    .A2(_1245_),
    .B(_1227_),
    .C(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5856_ (.I(\as2650.halted ),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5857_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5858_ (.A1(_1061_),
    .A2(_1246_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5859_ (.A1(_4032_),
    .A2(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5860_ (.I(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5861_ (.I(_1255_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5862_ (.I(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5863_ (.I(_0938_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5864_ (.I(_1219_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5865_ (.I(_1259_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5866_ (.I(_1049_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5867_ (.A1(_1215_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5868_ (.I(_1262_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5869_ (.A1(_1258_),
    .A2(_1260_),
    .B(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5870_ (.A1(_0872_),
    .A2(_1244_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5871_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5872_ (.A1(_1073_),
    .A2(_4300_),
    .A3(_4071_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5873_ (.A1(_4073_),
    .A2(_4077_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5874_ (.A1(_1267_),
    .A2(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5875_ (.A1(_1269_),
    .A2(_1222_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5876_ (.I(_1069_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5877_ (.I(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5878_ (.I(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5879_ (.A1(_1249_),
    .A2(_1266_),
    .B(_1270_),
    .C(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5880_ (.I(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5881_ (.A1(_1252_),
    .A2(_1257_),
    .A3(_1264_),
    .A4(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5882_ (.A1(_1228_),
    .A2(_1239_),
    .A3(_1250_),
    .A4(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5883_ (.I(_1225_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5884_ (.I(_1278_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5885_ (.A1(_0589_),
    .A2(_4308_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5886_ (.I(_0604_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5887_ (.I(_1281_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5888_ (.I(_1282_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5889_ (.I(_4109_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5890_ (.I(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5891_ (.I(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5892_ (.I(_1281_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5893_ (.A1(_4310_),
    .A2(_1245_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5894_ (.A1(_1287_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5895_ (.A1(\as2650.psu[5] ),
    .A2(_1283_),
    .B(_1286_),
    .C(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5896_ (.A1(_1280_),
    .A2(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5897_ (.A1(_1279_),
    .A2(_1291_),
    .B(_1277_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5898_ (.I(_0940_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5899_ (.I(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5900_ (.I(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5901_ (.A1(_1213_),
    .A2(_1277_),
    .B(_1292_),
    .C(_1295_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5902_ (.I(_0911_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5903_ (.I(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5904_ (.I(_1297_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5905_ (.A1(_1044_),
    .A2(_1298_),
    .A3(_1084_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5906_ (.I(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5907_ (.I(_1300_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5908_ (.I(_1300_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5909_ (.A1(\as2650.stack[0][8] ),
    .A2(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5910_ (.A1(_1190_),
    .A2(_1301_),
    .B(_1303_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5911_ (.I(_1299_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5912_ (.A1(\as2650.stack[0][9] ),
    .A2(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5913_ (.A1(_1200_),
    .A2(_1301_),
    .B(_1305_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5914_ (.A1(\as2650.stack[0][10] ),
    .A2(_1304_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5915_ (.A1(_1203_),
    .A2(_1301_),
    .B(_1306_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5916_ (.A1(\as2650.stack[0][11] ),
    .A2(_1304_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5917_ (.A1(_1205_),
    .A2(_1301_),
    .B(_1307_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5918_ (.A1(\as2650.stack[0][12] ),
    .A2(_1304_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5919_ (.A1(_1207_),
    .A2(_1302_),
    .B(_1308_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5920_ (.A1(\as2650.stack[0][13] ),
    .A2(_1300_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5921_ (.A1(_1209_),
    .A2(_1302_),
    .B(_1309_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5922_ (.A1(\as2650.stack[0][14] ),
    .A2(_1300_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5923_ (.A1(_1211_),
    .A2(_1302_),
    .B(_1310_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5924_ (.A1(_0804_),
    .A2(_0815_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5925_ (.A1(_4186_),
    .A2(_4355_),
    .A3(_0316_),
    .A4(_0412_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5926_ (.A1(_0700_),
    .A2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5927_ (.A1(_0511_),
    .A2(_0650_),
    .A3(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5928_ (.A1(_0800_),
    .A2(_0801_),
    .B(_0682_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5929_ (.A1(_0501_),
    .A2(_0627_),
    .A3(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5930_ (.I(_4293_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5931_ (.A1(_1317_),
    .A2(_4337_),
    .A3(_0298_),
    .A4(_0386_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5932_ (.A1(_4159_),
    .A2(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5933_ (.A1(_0388_),
    .A2(_0303_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5934_ (.A1(_4329_),
    .A2(_0305_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5935_ (.A1(_4156_),
    .A2(_4169_),
    .B(_4344_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5936_ (.A1(_1321_),
    .A2(_1322_),
    .B(_0386_),
    .C(_0298_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5937_ (.A1(_0384_),
    .A2(_1320_),
    .B1(_0496_),
    .B2(_0497_),
    .C(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5938_ (.A1(_0647_),
    .A2(_0639_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5939_ (.A1(_0625_),
    .A2(_0629_),
    .B(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5940_ (.A1(_1315_),
    .A2(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5941_ (.A1(_0800_),
    .A2(_0811_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5942_ (.A1(_1324_),
    .A2(_1316_),
    .B(_1327_),
    .C(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5943_ (.A1(_0698_),
    .A2(_0692_),
    .A3(_0802_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5944_ (.A1(\as2650.psl[1] ),
    .A2(_0803_),
    .B(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5945_ (.A1(_1329_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5946_ (.A1(\as2650.psl[1] ),
    .A2(_0803_),
    .A3(_1328_),
    .B(_4396_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5947_ (.I(_1091_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5948_ (.I(_1334_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5949_ (.I(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5950_ (.A1(_1332_),
    .A2(_1333_),
    .B(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5951_ (.A1(_1316_),
    .A2(_1319_),
    .B(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5952_ (.A1(_4396_),
    .A2(_1311_),
    .A3(_1314_),
    .B(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5953_ (.I(_4223_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5954_ (.I(_4087_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5955_ (.I(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5956_ (.I(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5957_ (.I(_4143_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5958_ (.A1(_4142_),
    .A2(_1343_),
    .A3(_1243_),
    .A4(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5959_ (.I(_1345_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5960_ (.A1(_1340_),
    .A2(_0778_),
    .A3(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5961_ (.I(_4294_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5962_ (.A1(_0333_),
    .A2(_4376_),
    .A3(_4188_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5963_ (.A1(_0711_),
    .A2(_0589_),
    .A3(_0517_),
    .A4(_0414_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5964_ (.A1(_1348_),
    .A2(_1349_),
    .A3(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5965_ (.I(_4037_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5966_ (.I(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5967_ (.I(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5968_ (.I(_1354_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5969_ (.A1(_1039_),
    .A2(_1346_),
    .B(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5970_ (.A1(_1351_),
    .A2(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5971_ (.I(_4362_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5972_ (.I(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5973_ (.I(_1359_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5974_ (.A1(_1347_),
    .A2(_1357_),
    .B(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5975_ (.I(_1359_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5976_ (.I(_4101_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5977_ (.I(_4224_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5978_ (.I(_1268_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5979_ (.A1(_1365_),
    .A2(_0602_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5980_ (.A1(_1364_),
    .A2(_0705_),
    .B(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5981_ (.A1(_1240_),
    .A2(_1241_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5982_ (.A1(_4164_),
    .A2(_4099_),
    .A3(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5983_ (.I(_1369_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5984_ (.I(_0723_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5985_ (.I(_1371_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5986_ (.I(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5987_ (.I(_1373_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5988_ (.I(\as2650.psl[6] ),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5989_ (.A1(_1375_),
    .A2(_1374_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5990_ (.A1(_0521_),
    .A2(_1374_),
    .B(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5991_ (.A1(_4007_),
    .A2(_1370_),
    .A3(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5992_ (.A1(_1349_),
    .A2(_1350_),
    .B(_0792_),
    .C(_1259_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5993_ (.A1(_0711_),
    .A2(_1260_),
    .B(_1379_),
    .C(_0938_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5994_ (.I(_1365_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5995_ (.A1(_1285_),
    .A2(_1378_),
    .B(_1380_),
    .C(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5996_ (.I(_4072_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5997_ (.A1(_1367_),
    .A2(_1382_),
    .B(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5998_ (.I(_1267_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5999_ (.I(_0602_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_0304_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6001_ (.I(_0346_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6002_ (.A1(_1387_),
    .A2(_0717_),
    .A3(_4390_),
    .A4(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6003_ (.A1(_0428_),
    .A2(_0714_),
    .A3(_1386_),
    .A4(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6004_ (.A1(_1385_),
    .A2(_0782_),
    .A3(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6005_ (.A1(_1363_),
    .A2(_1384_),
    .A3(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6006_ (.I(_0785_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6007_ (.A1(_1344_),
    .A2(_1222_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6008_ (.I(_1394_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6009_ (.I(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6010_ (.A1(_1393_),
    .A2(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6011_ (.I(_4243_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6012_ (.I(_1398_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6013_ (.I(_4392_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6014_ (.I(_1400_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6015_ (.I(net7),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6016_ (.I(_1402_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6017_ (.I(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6018_ (.I(_1404_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6019_ (.I(_0431_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6020_ (.I(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6021_ (.A1(_1399_),
    .A2(_1401_),
    .A3(_1405_),
    .A4(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6022_ (.I(_0540_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6023_ (.I(_1409_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6024_ (.I(_1410_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6025_ (.I(_1374_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6026_ (.A1(_1411_),
    .A2(_1287_),
    .A3(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6027_ (.A1(_1396_),
    .A2(_1408_),
    .A3(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6028_ (.A1(_1362_),
    .A2(_1392_),
    .A3(_1397_),
    .A4(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6029_ (.A1(_1217_),
    .A2(_1259_),
    .A3(_1262_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6030_ (.I(_4040_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6031_ (.A1(_1417_),
    .A2(_1341_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6032_ (.A1(_4145_),
    .A2(_0927_),
    .A3(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6033_ (.A1(_4292_),
    .A2(_1227_),
    .A3(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6034_ (.I(_4049_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6035_ (.I(_1269_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6036_ (.A1(_4080_),
    .A2(_1229_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6037_ (.A1(_1255_),
    .A2(_1422_),
    .A3(_1223_),
    .A4(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6038_ (.A1(_1421_),
    .A2(_1424_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6039_ (.A1(_4260_),
    .A2(_4291_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6040_ (.I(_4031_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6041_ (.A1(_1427_),
    .A2(_1247_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6042_ (.A1(_1428_),
    .A2(_4125_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6043_ (.I(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6044_ (.A1(_1426_),
    .A2(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6045_ (.A1(_1416_),
    .A2(_1420_),
    .B(_1425_),
    .C(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6046_ (.I(_4084_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6047_ (.A1(_1433_),
    .A2(_1394_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6048_ (.A1(_4007_),
    .A2(_1284_),
    .A3(_1217_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6049_ (.A1(_1341_),
    .A2(_4296_),
    .A3(_4331_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6050_ (.A1(_4038_),
    .A2(_1436_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6051_ (.A1(_1246_),
    .A2(_1247_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6052_ (.A1(_4102_),
    .A2(_1438_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6053_ (.I(_1439_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6054_ (.A1(_4007_),
    .A2(_1440_),
    .A3(_1245_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6055_ (.I(_1075_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6056_ (.I(_4105_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6057_ (.A1(_4361_),
    .A2(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6058_ (.A1(_1251_),
    .A2(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6059_ (.A1(_1442_),
    .A2(_1263_),
    .A3(_1278_),
    .A4(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6060_ (.A1(_1435_),
    .A2(_1437_),
    .A3(_1441_),
    .A4(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6061_ (.A1(_1434_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6062_ (.I(_1418_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6063_ (.I(_1342_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6064_ (.I(_4083_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6065_ (.A1(_1451_),
    .A2(_4193_),
    .A3(_1436_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6066_ (.A1(_4310_),
    .A2(_4116_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6067_ (.A1(_1450_),
    .A2(_1452_),
    .A3(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6068_ (.I(_1454_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _6069_ (.A1(_0405_),
    .A2(_1250_),
    .A3(_1449_),
    .B1(_1455_),
    .B2(_1345_),
    .B3(_4196_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6070_ (.A1(_1343_),
    .A2(_1091_),
    .A3(_4202_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6071_ (.A1(_4109_),
    .A2(_4225_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6072_ (.I(_1344_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6073_ (.I(_4100_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6074_ (.A1(_1242_),
    .A2(_1459_),
    .A3(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6075_ (.A1(_4260_),
    .A2(_4108_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6076_ (.A1(_4101_),
    .A2(_1418_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6077_ (.I(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6078_ (.A1(_4037_),
    .A2(_1453_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6079_ (.A1(_0640_),
    .A2(_1462_),
    .B1(_1464_),
    .B2(_1254_),
    .C(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6080_ (.A1(_1457_),
    .A2(_1458_),
    .A3(_1461_),
    .A4(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6081_ (.A1(_1432_),
    .A2(_1448_),
    .A3(_1456_),
    .A4(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6082_ (.A1(_1415_),
    .A2(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6083_ (.A1(_1339_),
    .A2(_1361_),
    .B(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6084_ (.I(_4285_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6085_ (.A1(_1375_),
    .A2(_1468_),
    .B(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6086_ (.A1(_1470_),
    .A2(_1472_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6087_ (.I(_1358_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6088_ (.I(_1473_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6089_ (.A1(_0804_),
    .A2(_0815_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6090_ (.A1(_4127_),
    .A2(_1475_),
    .B(_1337_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6091_ (.A1(_1340_),
    .A2(_1346_),
    .B(_1356_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6092_ (.A1(_1362_),
    .A2(_1397_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6093_ (.I(_4072_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6094_ (.A1(_1479_),
    .A2(_0782_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6095_ (.I(_1214_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6096_ (.A1(_1224_),
    .A2(_1417_),
    .A3(_4128_),
    .A4(_4335_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6097_ (.A1(_4006_),
    .A2(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6098_ (.I(_0430_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6099_ (.I(\as2650.psu[3] ),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6100_ (.A1(_0910_),
    .A2(_1403_),
    .B1(_1484_),
    .B2(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6101_ (.I(\as2650.psu[7] ),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6102_ (.I(_0783_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6103_ (.A1(_1487_),
    .A2(_1488_),
    .B1(_0605_),
    .B2(_1213_),
    .C1(_4393_),
    .C2(_0897_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6104_ (.I(\as2650.psu[4] ),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6105_ (.I(_1371_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6106_ (.I(net27),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6107_ (.A1(_1490_),
    .A2(_0540_),
    .B1(_1491_),
    .B2(_1492_),
    .C1(_0895_),
    .C2(_4242_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6108_ (.A1(_1486_),
    .A2(_1489_),
    .A3(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6109_ (.I(_0400_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6110_ (.I(net5),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6111_ (.A1(_1496_),
    .A2(_4249_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6112_ (.A1(_1484_),
    .A2(_1495_),
    .B1(_0536_),
    .B2(_0605_),
    .C(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6113_ (.I(net3),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6114_ (.I(_0527_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6115_ (.A1(_1499_),
    .A2(_0716_),
    .B1(_1482_),
    .B2(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6116_ (.I(net6),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6117_ (.A1(_0540_),
    .A2(_0427_),
    .B1(_0601_),
    .B2(_1372_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6118_ (.A1(_1502_),
    .A2(_1387_),
    .B1(_4389_),
    .B2(_0348_),
    .C(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6119_ (.A1(_1501_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6120_ (.I(\as2650.overflow ),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6121_ (.I(\as2650.psl[5] ),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6122_ (.A1(_1506_),
    .A2(_1403_),
    .B1(_0604_),
    .B2(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6123_ (.A1(\as2650.psl[7] ),
    .A2(_1499_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6124_ (.A1(_4173_),
    .A2(_4241_),
    .B1(_0430_),
    .B2(_4207_),
    .C(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6125_ (.I(\as2650.psl[1] ),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6126_ (.A1(_1375_),
    .A2(_0725_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6127_ (.A1(_1511_),
    .A2(_4392_),
    .B1(_0539_),
    .B2(_4015_),
    .C(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6128_ (.A1(_1508_),
    .A2(_1510_),
    .A3(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6129_ (.A1(_4005_),
    .A2(_1514_),
    .B(_1482_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6130_ (.A1(_1498_),
    .A2(_1505_),
    .B(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6131_ (.A1(_1232_),
    .A2(_1369_),
    .B1(_1483_),
    .B2(_1494_),
    .C(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6132_ (.I(\as2650.psl[7] ),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6133_ (.I(_1488_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6134_ (.I(_1076_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6135_ (.A1(_1518_),
    .A2(_1519_),
    .A3(_1520_),
    .A4(_1244_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6136_ (.A1(_1265_),
    .A2(_1517_),
    .A3(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6137_ (.I(_1499_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6138_ (.A1(_1518_),
    .A2(_1523_),
    .A3(_1266_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6139_ (.A1(_1522_),
    .A2(_1524_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6140_ (.A1(_0792_),
    .A2(_4294_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6141_ (.I(_4078_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6142_ (.I(_1527_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6143_ (.A1(_1481_),
    .A2(_1525_),
    .B(_1526_),
    .C(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6144_ (.A1(_1383_),
    .A2(_1366_),
    .A3(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6145_ (.A1(_1480_),
    .A2(_1530_),
    .B(_1396_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6146_ (.A1(_1474_),
    .A2(_1476_),
    .A3(_1477_),
    .B1(_1478_),
    .B2(_1531_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6147_ (.A1(_1518_),
    .A2(_1468_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6148_ (.A1(_1468_),
    .A2(_1532_),
    .B(_1533_),
    .C(_1295_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6149_ (.I(\as2650.r123_2[3][0] ),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(_1534_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6151_ (.I(\as2650.r123_2[3][1] ),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6152_ (.I(_1535_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6153_ (.I(\as2650.r123_2[3][2] ),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6154_ (.I(_1536_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6155_ (.I(\as2650.r123_2[3][3] ),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6156_ (.I(_1537_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6157_ (.I(\as2650.r123_2[3][4] ),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6158_ (.I(_1538_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6159_ (.I(\as2650.r123_2[3][5] ),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6160_ (.I(_1539_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6161_ (.I(\as2650.r123_2[3][6] ),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6162_ (.I(_1540_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6163_ (.I(\as2650.r123_2[3][7] ),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6164_ (.I(_1541_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6165_ (.I(_4006_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6166_ (.A1(_1427_),
    .A2(_4054_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6167_ (.I(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6168_ (.A1(_4073_),
    .A2(_1070_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6169_ (.I(_1545_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6170_ (.I(_1546_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6171_ (.I(_1547_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6172_ (.I(_1548_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6173_ (.I(_4035_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6174_ (.I(_4288_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6175_ (.I(_1427_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6176_ (.I(_4105_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6177_ (.A1(_0784_),
    .A2(_1553_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6178_ (.A1(_1550_),
    .A2(_1551_),
    .A3(_1552_),
    .A4(_1554_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6179_ (.A1(_1544_),
    .A2(_1549_),
    .B(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6180_ (.I(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6181_ (.A1(_1542_),
    .A2(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6182_ (.I(_1399_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6183_ (.I(_1057_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6184_ (.A1(_4032_),
    .A2(_1427_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6185_ (.I(_1561_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6186_ (.A1(_1560_),
    .A2(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6187_ (.A1(_1551_),
    .A2(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6188_ (.I(_1564_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6189_ (.A1(_1559_),
    .A2(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6190_ (.I(_4044_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6191_ (.I(_1567_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6192_ (.I(_1568_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6193_ (.A1(_1569_),
    .A2(_1563_),
    .A3(_1555_),
    .A4(_1549_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6194_ (.A1(_1558_),
    .A2(_1566_),
    .A3(_1570_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6195_ (.A1(_0945_),
    .A2(_1557_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6196_ (.I(_1401_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6197_ (.I(_1564_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6198_ (.A1(_1572_),
    .A2(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6199_ (.A1(_1570_),
    .A2(_1571_),
    .A3(_1574_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6200_ (.I(_0349_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6201_ (.I(_1565_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6202_ (.I(_1224_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6203_ (.I(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6204_ (.A1(_1578_),
    .A2(_1565_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6205_ (.A1(_1575_),
    .A2(_1576_),
    .B(_1579_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6206_ (.I(_1442_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6207_ (.A1(_1580_),
    .A2(_1544_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6208_ (.A1(_1231_),
    .A2(_1555_),
    .A3(_1549_),
    .A4(_1581_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6209_ (.A1(_1283_),
    .A2(_1565_),
    .B1(_1556_),
    .B2(_1231_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6210_ (.A1(_1582_),
    .A2(_1583_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6211_ (.I(_1412_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6212_ (.A1(_1584_),
    .A2(_1576_),
    .B1(_1557_),
    .B2(_1243_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6213_ (.I(_1585_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6214_ (.I(_1393_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6215_ (.A1(_1586_),
    .A2(_1573_),
    .B1(_1557_),
    .B2(_1459_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6216_ (.I(_1587_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6217_ (.I(_4188_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6218_ (.I(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6219_ (.I(_1589_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6220_ (.A1(_0861_),
    .A2(_1093_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6221_ (.I(_1591_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6222_ (.A1(_1592_),
    .A2(_1160_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6223_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6224_ (.I(_1594_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6225_ (.I(\as2650.pc[0] ),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6226_ (.I(_1596_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6227_ (.I(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6228_ (.I(_1598_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6229_ (.A1(_1067_),
    .A2(_1068_),
    .A3(_1071_),
    .B(_1080_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6230_ (.A1(_0861_),
    .A2(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6231_ (.I(_1601_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6232_ (.A1(_1602_),
    .A2(_1147_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6233_ (.I(_1603_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6234_ (.I(_1082_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6235_ (.A1(_1044_),
    .A2(_0971_),
    .A3(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6236_ (.I(_1606_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6237_ (.I(_1593_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6238_ (.A1(_1599_),
    .A2(_1604_),
    .B1(_1607_),
    .B2(\as2650.stack[5][0] ),
    .C(_1608_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6239_ (.A1(_1590_),
    .A2(_1595_),
    .B(_1609_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6240_ (.I(_4230_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6241_ (.I(_1610_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6242_ (.I(\as2650.pc[1] ),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6243_ (.I(_1612_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6244_ (.I(_1613_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6245_ (.I(_1614_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6246_ (.I(_1606_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6247_ (.A1(\as2650.stack[5][1] ),
    .A2(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6248_ (.A1(_1615_),
    .A2(_1604_),
    .B(_1594_),
    .C(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6249_ (.A1(_1611_),
    .A2(_1595_),
    .B(_1618_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6250_ (.I(_0981_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6251_ (.I(_1619_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6252_ (.I(\as2650.pc[2] ),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6253_ (.I(_1621_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6254_ (.I(_1622_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6255_ (.I(_1623_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6256_ (.I(_1603_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6257_ (.A1(_1624_),
    .A2(_1625_),
    .B1(_1607_),
    .B2(\as2650.stack[5][2] ),
    .C(_1608_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6258_ (.A1(_1620_),
    .A2(_1595_),
    .B(_1626_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6259_ (.I(_0415_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6260_ (.I(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6261_ (.I(_1628_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6262_ (.I(\as2650.pc[3] ),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6263_ (.I(_1630_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6264_ (.I(_1631_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6265_ (.A1(\as2650.stack[5][3] ),
    .A2(_1616_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6266_ (.A1(_1632_),
    .A2(_1604_),
    .B(_1594_),
    .C(_1633_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6267_ (.A1(_1629_),
    .A2(_1595_),
    .B(_1634_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6268_ (.I(_0518_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6269_ (.I(_1635_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6270_ (.I(_1594_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6271_ (.I(\as2650.pc[4] ),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6272_ (.I(_1638_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6273_ (.I(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6274_ (.A1(_1640_),
    .A2(_1625_),
    .B1(_1607_),
    .B2(\as2650.stack[5][4] ),
    .C(_1608_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6275_ (.A1(_1636_),
    .A2(_1637_),
    .B(_1641_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6276_ (.I(_0590_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6277_ (.I(\as2650.pc[5] ),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6278_ (.I(_1643_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6279_ (.I(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6280_ (.I(_1645_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6281_ (.A1(_1646_),
    .A2(_1625_),
    .B1(_1607_),
    .B2(\as2650.stack[5][5] ),
    .C(_1593_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6282_ (.A1(_1642_),
    .A2(_1637_),
    .B(_1647_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6283_ (.I(_0713_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6284_ (.I(_1648_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6285_ (.I(\as2650.pc[6] ),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6286_ (.I(_1650_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6287_ (.A1(_1651_),
    .A2(_1625_),
    .B1(_1616_),
    .B2(\as2650.stack[5][6] ),
    .C(_1593_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6288_ (.A1(_1649_),
    .A2(_1637_),
    .B(_1652_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6289_ (.I(_1040_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6290_ (.I(_1653_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6291_ (.I(\as2650.pc[7] ),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6292_ (.I(_1655_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6293_ (.I(_1656_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6294_ (.A1(\as2650.stack[5][7] ),
    .A2(_1616_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6295_ (.A1(_1657_),
    .A2(_1604_),
    .B(_1608_),
    .C(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6296_ (.A1(_1654_),
    .A2(_1637_),
    .B(_1659_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6297_ (.A1(_1592_),
    .A2(_1147_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6298_ (.I(_1660_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6299_ (.I(_1661_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6300_ (.A1(_0910_),
    .A2(_1296_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6301_ (.A1(_1663_),
    .A2(_1605_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6302_ (.I(_1664_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6303_ (.I(_1596_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6304_ (.I(_1666_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6305_ (.A1(_1667_),
    .A2(_1665_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6306_ (.A1(\as2650.stack[4][0] ),
    .A2(_1665_),
    .B(_1668_),
    .C(_1661_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6307_ (.A1(_1590_),
    .A2(_1662_),
    .B(_1669_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6308_ (.I(_1614_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6309_ (.A1(_0967_),
    .A2(_1602_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6310_ (.I(_1664_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6311_ (.A1(\as2650.stack[4][1] ),
    .A2(_1672_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6312_ (.A1(_1670_),
    .A2(_1671_),
    .B(_1673_),
    .C(_1661_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6313_ (.A1(_1611_),
    .A2(_1662_),
    .B(_1674_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6314_ (.I(_1619_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6315_ (.I(_1661_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6316_ (.I(_1672_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6317_ (.A1(\as2650.stack[4][2] ),
    .A2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6318_ (.I(_1623_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6319_ (.I(_1671_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6320_ (.I(_1660_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6321_ (.A1(_1679_),
    .A2(_1680_),
    .B(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6322_ (.A1(_1675_),
    .A2(_1676_),
    .B1(_1678_),
    .B2(_1682_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6323_ (.I(\as2650.pc[3] ),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6324_ (.I(_1683_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6325_ (.A1(_1684_),
    .A2(_1672_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6326_ (.A1(\as2650.stack[4][3] ),
    .A2(_1665_),
    .B(_1685_),
    .C(_1660_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6327_ (.A1(_1629_),
    .A2(_1662_),
    .B(_1686_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6328_ (.I(\as2650.pc[4] ),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6329_ (.I(_1687_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6330_ (.I(_1688_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6331_ (.A1(_1689_),
    .A2(_1672_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6332_ (.A1(\as2650.stack[4][4] ),
    .A2(_1665_),
    .B(_1690_),
    .C(_1660_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6333_ (.A1(_1636_),
    .A2(_1662_),
    .B(_1691_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6334_ (.A1(\as2650.stack[4][5] ),
    .A2(_1677_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6335_ (.I(_1645_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6336_ (.A1(_1693_),
    .A2(_1680_),
    .B(_1681_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6337_ (.A1(_1642_),
    .A2(_1676_),
    .B1(_1692_),
    .B2(_1694_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6338_ (.A1(\as2650.stack[4][6] ),
    .A2(_1677_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6339_ (.I(_1651_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6340_ (.A1(_1696_),
    .A2(_1680_),
    .B(_1681_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6341_ (.A1(_1648_),
    .A2(_1676_),
    .B1(_1695_),
    .B2(_1697_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6342_ (.I(_1653_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6343_ (.A1(\as2650.stack[4][7] ),
    .A2(_1677_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6344_ (.A1(_1657_),
    .A2(_1680_),
    .B(_1681_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6345_ (.A1(_1698_),
    .A2(_1676_),
    .B1(_1699_),
    .B2(_1700_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6346_ (.I(\as2650.r123[3][0] ),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6347_ (.I(_1701_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6348_ (.I(\as2650.r123[3][1] ),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6349_ (.I(_1702_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6350_ (.I(\as2650.r123[3][2] ),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6351_ (.I(_1703_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6352_ (.I(\as2650.r123[3][3] ),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6353_ (.I(_1704_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6354_ (.I(\as2650.r123[3][4] ),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6355_ (.I(_1705_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6356_ (.I(\as2650.r123[3][5] ),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6357_ (.I(_1706_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6358_ (.I(\as2650.r123[3][6] ),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6359_ (.I(_1707_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6360_ (.I(\as2650.r123[3][7] ),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6361_ (.I(_1708_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6362_ (.I(_1589_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6363_ (.A1(_0967_),
    .A2(_1592_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6364_ (.I(_1710_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6365_ (.I(_1711_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6366_ (.I(_0910_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6367_ (.A1(_1713_),
    .A2(_0969_),
    .A3(_1605_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6368_ (.I(_1714_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6369_ (.A1(\as2650.stack[3][0] ),
    .A2(_1715_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6370_ (.A1(_1174_),
    .A2(_1048_),
    .A3(_1601_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6371_ (.I(_1717_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6372_ (.I(_1710_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6373_ (.A1(_1599_),
    .A2(_1718_),
    .B(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6374_ (.A1(_1709_),
    .A2(_1712_),
    .B1(_1716_),
    .B2(_1720_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6375_ (.I(_1610_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6376_ (.I(_1711_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6377_ (.A1(\as2650.stack[3][1] ),
    .A2(_1715_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6378_ (.A1(_1615_),
    .A2(_1718_),
    .B(_1719_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6379_ (.A1(_1721_),
    .A2(_1722_),
    .B1(_1723_),
    .B2(_1724_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6380_ (.A1(\as2650.stack[3][2] ),
    .A2(_1715_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6381_ (.A1(_1679_),
    .A2(_1718_),
    .B(_1719_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6382_ (.A1(_1675_),
    .A2(_1722_),
    .B1(_1725_),
    .B2(_1726_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6383_ (.I(_1628_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6384_ (.A1(\as2650.stack[3][3] ),
    .A2(_1715_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6385_ (.I(_1632_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6386_ (.A1(_1729_),
    .A2(_1718_),
    .B(_1719_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6387_ (.A1(_1727_),
    .A2(_1722_),
    .B1(_1728_),
    .B2(_1730_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6388_ (.I(_1714_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6389_ (.A1(_1689_),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6390_ (.A1(\as2650.stack[3][4] ),
    .A2(_1731_),
    .B(_1732_),
    .C(_1711_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6391_ (.A1(_1636_),
    .A2(_1712_),
    .B(_1733_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6392_ (.I(_0590_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6393_ (.A1(\as2650.stack[3][5] ),
    .A2(_1731_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6394_ (.A1(_1693_),
    .A2(_1717_),
    .B(_1711_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6395_ (.A1(_1734_),
    .A2(_1722_),
    .B1(_1735_),
    .B2(_1736_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6396_ (.I(\as2650.pc[6] ),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6397_ (.I(_1737_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6398_ (.A1(_1738_),
    .A2(_1714_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6399_ (.A1(\as2650.stack[3][6] ),
    .A2(_1731_),
    .B(_1739_),
    .C(_1710_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6400_ (.A1(_1649_),
    .A2(_1712_),
    .B(_1740_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6401_ (.I(_1656_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6402_ (.A1(\as2650.stack[3][7] ),
    .A2(_1714_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6403_ (.A1(_1741_),
    .A2(_1717_),
    .B(_1710_),
    .C(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6404_ (.A1(_1654_),
    .A2(_1712_),
    .B(_1743_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6405_ (.A1(_1174_),
    .A2(_1048_),
    .A3(_1591_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6406_ (.I(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6407_ (.I(_1745_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6408_ (.I(_1173_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6409_ (.A1(_1747_),
    .A2(_1177_),
    .A3(_1601_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6410_ (.I(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6411_ (.I(_1082_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6412_ (.A1(_1713_),
    .A2(_0973_),
    .A3(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6413_ (.I(_1751_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6414_ (.A1(_1599_),
    .A2(_1749_),
    .B1(_1752_),
    .B2(\as2650.stack[2][0] ),
    .C(_1745_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6415_ (.A1(_1590_),
    .A2(_1746_),
    .B(_1753_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6416_ (.A1(_1670_),
    .A2(_1749_),
    .B1(_1752_),
    .B2(\as2650.stack[2][1] ),
    .C(_1745_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6417_ (.A1(_1611_),
    .A2(_1746_),
    .B(_1754_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6418_ (.I(_1744_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6419_ (.A1(_1624_),
    .A2(_1749_),
    .B1(_1752_),
    .B2(\as2650.stack[2][2] ),
    .C(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6420_ (.A1(_1620_),
    .A2(_1746_),
    .B(_1756_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6421_ (.A1(_1632_),
    .A2(_1749_),
    .B1(_1752_),
    .B2(\as2650.stack[2][3] ),
    .C(_1755_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6422_ (.A1(_1629_),
    .A2(_1746_),
    .B(_1757_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6423_ (.I(_1745_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6424_ (.I(_1748_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6425_ (.I(_1751_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6426_ (.A1(_1639_),
    .A2(_1759_),
    .B1(_1760_),
    .B2(\as2650.stack[2][4] ),
    .C(_1755_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6427_ (.A1(_1636_),
    .A2(_1758_),
    .B(_1761_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6428_ (.A1(_1646_),
    .A2(_1759_),
    .B1(_1760_),
    .B2(\as2650.stack[2][5] ),
    .C(_1755_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6429_ (.A1(_1642_),
    .A2(_1758_),
    .B(_1762_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6430_ (.A1(_1651_),
    .A2(_1759_),
    .B1(_1760_),
    .B2(\as2650.stack[2][6] ),
    .C(_1744_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6431_ (.A1(_1649_),
    .A2(_1758_),
    .B(_1763_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6432_ (.A1(_1741_),
    .A2(_1759_),
    .B1(_1760_),
    .B2(\as2650.stack[2][7] ),
    .C(_1744_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6433_ (.A1(_1654_),
    .A2(_1758_),
    .B(_1764_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6434_ (.I(_1667_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6435_ (.A1(_1043_),
    .A2(_1194_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6436_ (.A1(_1082_),
    .A2(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6437_ (.I(_1767_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6438_ (.I(_1767_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6439_ (.A1(\as2650.stack[1][0] ),
    .A2(_1769_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6440_ (.A1(_1765_),
    .A2(_1768_),
    .B(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6441_ (.A1(_1146_),
    .A2(_1177_),
    .A3(_1591_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6442_ (.I(_1772_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6443_ (.I(_1773_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6444_ (.I0(_1771_),
    .I1(_4306_),
    .S(_1774_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6445_ (.I(_1775_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6446_ (.I0(_1614_),
    .I1(\as2650.stack[1][1] ),
    .S(_1769_),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6447_ (.I(_4377_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6448_ (.I(_1772_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6449_ (.I0(_1776_),
    .I1(_1777_),
    .S(_1778_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6450_ (.I(_1779_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6451_ (.A1(_1623_),
    .A2(_1750_),
    .A3(_1766_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6452_ (.A1(\as2650.stack[1][2] ),
    .A2(_1768_),
    .B(_1780_),
    .C(_1773_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6453_ (.A1(_1620_),
    .A2(_1774_),
    .B(_1781_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6454_ (.I(_1767_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6455_ (.A1(_1684_),
    .A2(_1782_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6456_ (.A1(\as2650.stack[1][3] ),
    .A2(_1768_),
    .B(_1783_),
    .C(_1773_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6457_ (.A1(_1629_),
    .A2(_1774_),
    .B(_1784_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6458_ (.A1(\as2650.stack[1][4] ),
    .A2(_1769_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6459_ (.A1(_1689_),
    .A2(_1782_),
    .B(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6460_ (.I0(_1786_),
    .I1(_1000_),
    .S(_1778_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6461_ (.I(_1787_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6462_ (.I0(_1645_),
    .I1(\as2650.stack[1][5] ),
    .S(_1767_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6463_ (.I0(_1788_),
    .I1(_1022_),
    .S(_1778_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6464_ (.I(_1789_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6465_ (.A1(\as2650.stack[1][6] ),
    .A2(_1769_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6466_ (.A1(_1738_),
    .A2(_1782_),
    .B(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6467_ (.I0(_1791_),
    .I1(_1028_),
    .S(_1778_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6468_ (.I(_1792_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6469_ (.I(_1655_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6470_ (.I(_1793_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6471_ (.A1(_1794_),
    .A2(_1782_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6472_ (.A1(\as2650.stack[1][7] ),
    .A2(_1768_),
    .B(_1795_),
    .C(_1773_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6473_ (.A1(_1654_),
    .A2(_1774_),
    .B(_1796_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6474_ (.I(_0937_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6475_ (.A1(_4286_),
    .A2(_4110_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6476_ (.I(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6477_ (.A1(_1797_),
    .A2(_4314_),
    .A3(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6478_ (.I(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6479_ (.A1(_0291_),
    .A2(_1095_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6480_ (.I(_1802_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6481_ (.A1(_4131_),
    .A2(_1798_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6482_ (.I(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6483_ (.I(_1805_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6484_ (.A1(_4366_),
    .A2(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6485_ (.I(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6486_ (.A1(_4098_),
    .A2(_1805_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6487_ (.I(_1809_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6488_ (.A1(_4310_),
    .A2(_1095_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6489_ (.A1(_4082_),
    .A2(_1811_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6490_ (.I(_1812_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6491_ (.A1(_4196_),
    .A2(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6492_ (.I(_1814_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6493_ (.I(_1815_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6494_ (.A1(_4202_),
    .A2(_1813_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6495_ (.I(_1817_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6496_ (.I(_1818_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6497_ (.A1(_4225_),
    .A2(_1812_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6498_ (.I(_1820_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6499_ (.A1(_0353_),
    .A2(_1804_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6500_ (.I(_1822_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6501_ (.A1(_1241_),
    .A2(_1394_),
    .A3(_1248_),
    .A4(_1804_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6502_ (.A1(_4250_),
    .A2(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6503_ (.A1(_4243_),
    .A2(_1823_),
    .B(_1825_),
    .C(_1820_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6504_ (.A1(_4239_),
    .A2(_1821_),
    .B(_1826_),
    .C(_1818_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6505_ (.A1(_4224_),
    .A2(_1819_),
    .B(_1827_),
    .C(_1815_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6506_ (.I(_1809_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6507_ (.A1(_1588_),
    .A2(_1816_),
    .B(_1828_),
    .C(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6508_ (.A1(_4272_),
    .A2(_1810_),
    .B(_1830_),
    .C(_1807_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6509_ (.I(_1802_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6510_ (.A1(_4279_),
    .A2(_1808_),
    .B(_1831_),
    .C(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6511_ (.A1(_4186_),
    .A2(_1803_),
    .B(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6512_ (.A1(_1801_),
    .A2(_1834_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6513_ (.I(_1820_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6514_ (.I(_1836_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6515_ (.I(_1817_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6516_ (.I(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6517_ (.A1(_4045_),
    .A2(_4061_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6518_ (.A1(_1840_),
    .A2(_1806_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6519_ (.I(_1814_),
    .Z(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6520_ (.I(_0865_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6521_ (.A1(_0864_),
    .A2(_1843_),
    .A3(_1805_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6522_ (.I(_1056_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6523_ (.A1(_4361_),
    .A2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6524_ (.A1(_0641_),
    .A2(_4127_),
    .A3(_4132_),
    .A4(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6525_ (.A1(_1847_),
    .A2(_1095_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6526_ (.A1(_1842_),
    .A2(_1824_),
    .A3(_1844_),
    .A4(_1848_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6527_ (.A1(_1837_),
    .A2(_1839_),
    .A3(_1841_),
    .A4(_1849_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6528_ (.A1(_1520_),
    .A2(_1850_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6529_ (.I(_1851_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6530_ (.I(_1822_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6531_ (.I(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6532_ (.I(_1854_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6533_ (.A1(_4133_),
    .A2(_1799_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6534_ (.A1(_0864_),
    .A2(_1843_),
    .A3(_1806_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6535_ (.A1(_1069_),
    .A2(_1269_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6536_ (.I(_1858_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6537_ (.A1(_1859_),
    .A2(_1813_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6538_ (.A1(_1816_),
    .A2(_1857_),
    .A3(_1841_),
    .A4(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6539_ (.A1(_1855_),
    .A2(_1856_),
    .A3(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6540_ (.A1(_1520_),
    .A2(_1862_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6541_ (.A1(_1801_),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6542_ (.I(_1864_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6543_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6544_ (.I(_1801_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6545_ (.A1(_0825_),
    .A2(_0855_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6546_ (.A1(_0820_),
    .A2(_0856_),
    .B(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6547_ (.A1(_0747_),
    .A2(_0829_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6548_ (.A1(_1870_),
    .A2(_0822_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6549_ (.A1(_0828_),
    .A2(_0854_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6550_ (.A1(_1871_),
    .A2(_0853_),
    .B(_1872_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6551_ (.A1(_4210_),
    .A2(_4321_),
    .A3(_0832_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6552_ (.A1(_0758_),
    .A2(_0837_),
    .A3(_0831_),
    .B(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6553_ (.A1(_0836_),
    .A2(_0852_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6554_ (.A1(_0836_),
    .A2(_0852_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6555_ (.A1(_0834_),
    .A2(_1876_),
    .B(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6556_ (.A1(_0837_),
    .A2(_0840_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6557_ (.A1(_0837_),
    .A2(_0840_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6558_ (.A1(_0838_),
    .A2(_1879_),
    .B(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6559_ (.A1(_4209_),
    .A2(_4416_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6560_ (.A1(_1881_),
    .A2(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6561_ (.A1(_0847_),
    .A2(_0850_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6562_ (.A1(_0841_),
    .A2(_0851_),
    .B(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6563_ (.A1(_0592_),
    .A2(_0369_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6564_ (.A1(_0751_),
    .A2(_0465_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6565_ (.A1(_4229_),
    .A2(_0839_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6566_ (.A1(_1887_),
    .A2(_1888_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6567_ (.A1(_1886_),
    .A2(_1889_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6568_ (.A1(_0563_),
    .A2(_0765_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6569_ (.A1(_4382_),
    .A2(_0526_),
    .B1(_0845_),
    .B2(_4375_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6570_ (.A1(_0762_),
    .A2(_1891_),
    .B1(_1892_),
    .B2(_0848_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6571_ (.A1(_0416_),
    .A2(_0560_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6572_ (.A1(_0335_),
    .A2(_0842_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6573_ (.A1(_1891_),
    .A2(_1894_),
    .A3(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6574_ (.A1(_1893_),
    .A2(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6575_ (.A1(_1890_),
    .A2(_1897_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6576_ (.A1(_1885_),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6577_ (.A1(_1883_),
    .A2(_1899_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6578_ (.A1(_1878_),
    .A2(_1900_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6579_ (.A1(_1875_),
    .A2(_1901_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6580_ (.A1(_1869_),
    .A2(_1873_),
    .A3(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6581_ (.A1(_1867_),
    .A2(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6582_ (.A1(_1835_),
    .A2(_1852_),
    .B(_1866_),
    .C(_1904_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6583_ (.I(_1800_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6584_ (.A1(_4061_),
    .A2(_1811_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6585_ (.I(_1906_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6586_ (.I(_1842_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6587_ (.I(_1818_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6588_ (.I(_1853_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6589_ (.A1(_4106_),
    .A2(_1805_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6590_ (.A1(_4400_),
    .A2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6591_ (.A1(_1400_),
    .A2(_1910_),
    .B(_1912_),
    .C(_1821_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6592_ (.A1(_0355_),
    .A2(_1837_),
    .B(_1838_),
    .C(_1913_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6593_ (.A1(_4379_),
    .A2(_1909_),
    .B(_1914_),
    .C(_1842_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6594_ (.A1(_4230_),
    .A2(_1908_),
    .B(_1829_),
    .C(_1915_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6595_ (.A1(_4263_),
    .A2(_1811_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6596_ (.I(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6597_ (.A1(_4374_),
    .A2(_1918_),
    .B(_1906_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6598_ (.A1(_4359_),
    .A2(_1907_),
    .B1(_1916_),
    .B2(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6599_ (.A1(_1848_),
    .A2(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6600_ (.A1(_4355_),
    .A2(_1803_),
    .B(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6601_ (.A1(_1905_),
    .A2(_1922_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6602_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_1865_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6603_ (.A1(_1873_),
    .A2(_1902_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6604_ (.A1(_1873_),
    .A2(_1902_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6605_ (.A1(_1869_),
    .A2(_1925_),
    .B(_1926_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6606_ (.A1(_1878_),
    .A2(_1900_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6607_ (.A1(_1875_),
    .A2(_1901_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6608_ (.A1(_1928_),
    .A2(_1929_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6609_ (.A1(_1881_),
    .A2(_1882_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6610_ (.A1(_1885_),
    .A2(_1898_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6611_ (.A1(_1883_),
    .A2(_1899_),
    .B(_1932_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6612_ (.A1(_4376_),
    .A2(_0470_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6613_ (.I(_0839_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6614_ (.I(_1935_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6615_ (.A1(_0588_),
    .A2(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6616_ (.A1(_1934_),
    .A2(_1937_),
    .B1(_1889_),
    .B2(_1886_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6617_ (.A1(_1893_),
    .A2(_1896_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6618_ (.A1(_1890_),
    .A2(_1897_),
    .B(_1939_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6619_ (.A1(_4208_),
    .A2(_0369_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6620_ (.A1(\as2650.r0[6] ),
    .A2(_4381_),
    .A3(_1935_),
    .A4(_0466_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6621_ (.A1(_4382_),
    .A2(_1935_),
    .B1(_0467_),
    .B2(_0592_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6622_ (.A1(_1942_),
    .A2(_1943_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6623_ (.A1(_1941_),
    .A2(_1944_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6624_ (.A1(\as2650.r0[3] ),
    .A2(_0765_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6625_ (.A1(_1891_),
    .A2(_1895_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6626_ (.A1(_0849_),
    .A2(_1946_),
    .B1(_1947_),
    .B2(_1894_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6627_ (.A1(_0416_),
    .A2(_0524_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6628_ (.A1(_1946_),
    .A2(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6629_ (.I(_0561_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6630_ (.A1(_0751_),
    .A2(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6631_ (.A1(_1950_),
    .A2(_1952_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6632_ (.A1(_1948_),
    .A2(_1953_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6633_ (.A1(_1945_),
    .A2(_1954_),
    .Z(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6634_ (.A1(_1940_),
    .A2(_1955_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6635_ (.A1(_1938_),
    .A2(_1956_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6636_ (.A1(_1933_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6637_ (.A1(_1931_),
    .A2(_1958_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6638_ (.A1(_1927_),
    .A2(_1930_),
    .A3(_1959_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6639_ (.A1(_1867_),
    .A2(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6640_ (.A1(_1852_),
    .A2(_1923_),
    .B(_1924_),
    .C(_1961_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6641_ (.I(_1851_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6642_ (.A1(_4294_),
    .A2(_4301_),
    .A3(_1096_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6643_ (.I(_1963_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6644_ (.I(_1856_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6645_ (.I(_1917_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6646_ (.A1(_0349_),
    .A2(_1855_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6647_ (.I(_1820_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6648_ (.A1(_0357_),
    .A2(_1855_),
    .B(_1967_),
    .C(_1968_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6649_ (.A1(_1495_),
    .A2(_1837_),
    .B(_1909_),
    .C(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6650_ (.I(_1815_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6651_ (.A1(_1387_),
    .A2(_1839_),
    .B(_1970_),
    .C(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6652_ (.A1(_0883_),
    .A2(_4116_),
    .A3(_1811_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6653_ (.A1(_0334_),
    .A2(_1973_),
    .B(_1918_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6654_ (.A1(_0331_),
    .A2(_1966_),
    .B1(_1972_),
    .B2(_1974_),
    .C(_1906_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6655_ (.A1(_0327_),
    .A2(_1907_),
    .B(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6656_ (.A1(_0316_),
    .A2(_1965_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6657_ (.A1(_1965_),
    .A2(_1976_),
    .B(_1977_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6658_ (.A1(_1964_),
    .A2(_1978_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6659_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_1865_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6660_ (.A1(_1941_),
    .A2(_1944_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6661_ (.A1(_1942_),
    .A2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6662_ (.A1(_1948_),
    .A2(_1953_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6663_ (.A1(_1945_),
    .A2(_1954_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6664_ (.A1(_1983_),
    .A2(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6665_ (.A1(_4208_),
    .A2(_1935_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6666_ (.A1(_0756_),
    .A2(_1986_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6667_ (.A1(_0337_),
    .A2(_1936_),
    .B1(_0470_),
    .B2(_4209_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6668_ (.A1(_1987_),
    .A2(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6669_ (.A1(_0417_),
    .A2(_0845_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6670_ (.A1(_1895_),
    .A2(_1990_),
    .B1(_1950_),
    .B2(_1952_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6671_ (.A1(_0751_),
    .A2(_0842_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6672_ (.A1(_1990_),
    .A2(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6673_ (.A1(_0593_),
    .A2(_1951_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6674_ (.A1(_1993_),
    .A2(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6675_ (.A1(_1991_),
    .A2(_1995_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6676_ (.A1(_1989_),
    .A2(_1996_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6677_ (.A1(_1985_),
    .A2(_1997_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6678_ (.A1(_1982_),
    .A2(_1998_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6679_ (.A1(_1940_),
    .A2(_1955_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6680_ (.A1(_1938_),
    .A2(_1956_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6681_ (.A1(_2000_),
    .A2(_2001_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6682_ (.A1(_1999_),
    .A2(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6683_ (.A1(_1933_),
    .A2(_1957_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6684_ (.A1(_1931_),
    .A2(_1958_),
    .B(_2004_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6685_ (.A1(_2003_),
    .A2(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6686_ (.A1(_1930_),
    .A2(_1959_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6687_ (.A1(_1930_),
    .A2(_1959_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6688_ (.A1(_1927_),
    .A2(_2007_),
    .B(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6689_ (.A1(_2006_),
    .A2(_2009_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6690_ (.A1(_1867_),
    .A2(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6691_ (.A1(_1962_),
    .A2(_1979_),
    .B(_1980_),
    .C(_2011_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6692_ (.I(_1963_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6693_ (.I(_2012_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6694_ (.I(_4390_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6695_ (.A1(_0436_),
    .A2(_1823_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6696_ (.A1(_0431_),
    .A2(_1910_),
    .B(_2015_),
    .C(_1821_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6697_ (.A1(_0427_),
    .A2(_1837_),
    .B(_1819_),
    .C(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6698_ (.A1(_2014_),
    .A2(_1839_),
    .B(_2017_),
    .C(_1816_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6699_ (.A1(_0414_),
    .A2(_1973_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6700_ (.A1(_2018_),
    .A2(_2019_),
    .B(_1918_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6701_ (.A1(_0452_),
    .A2(_1966_),
    .B(_1907_),
    .C(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6702_ (.A1(_0458_),
    .A2(_1808_),
    .B(_1802_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6703_ (.A1(_2021_),
    .A2(_2022_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6704_ (.A1(_0413_),
    .A2(_1965_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6705_ (.A1(_2023_),
    .A2(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6706_ (.A1(_2013_),
    .A2(_2025_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6707_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_1865_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6708_ (.A1(_2000_),
    .A2(_2001_),
    .B(_1999_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6709_ (.A1(_2003_),
    .A2(_2005_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6710_ (.A1(_2006_),
    .A2(_2009_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6711_ (.A1(_2029_),
    .A2(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6712_ (.A1(_1991_),
    .A2(_1995_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6713_ (.A1(_1989_),
    .A2(_1996_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6714_ (.A1(_2032_),
    .A2(_2033_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6715_ (.A1(_0418_),
    .A2(_1936_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6716_ (.I(_0845_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6717_ (.A1(_0533_),
    .A2(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6718_ (.A1(_1949_),
    .A2(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6719_ (.A1(_1993_),
    .A2(_1994_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6720_ (.A1(_2038_),
    .A2(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6721_ (.A1(_4208_),
    .A2(_1951_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6722_ (.A1(_0592_),
    .A2(_0842_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6723_ (.A1(_2037_),
    .A2(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6724_ (.A1(_2041_),
    .A2(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6725_ (.A1(_2040_),
    .A2(_2044_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6726_ (.A1(_2035_),
    .A2(_2045_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6727_ (.I(_2046_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6728_ (.A1(_2034_),
    .A2(_2047_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6729_ (.A1(_1987_),
    .A2(_2048_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6730_ (.A1(_1985_),
    .A2(_1997_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6731_ (.A1(_1942_),
    .A2(_1981_),
    .B(_1998_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6732_ (.A1(_2050_),
    .A2(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6733_ (.A1(_2049_),
    .A2(_2052_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6734_ (.A1(_2028_),
    .A2(_2031_),
    .A3(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6735_ (.A1(_1867_),
    .A2(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6736_ (.A1(_1962_),
    .A2(_2026_),
    .B(_2027_),
    .C(_2055_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6737_ (.I(_1807_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6738_ (.A1(_0543_),
    .A2(_1823_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6739_ (.A1(_1409_),
    .A2(_1910_),
    .B(_2057_),
    .C(_1836_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6740_ (.A1(_0537_),
    .A2(_1968_),
    .B(_1838_),
    .C(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6741_ (.A1(_1388_),
    .A2(_1909_),
    .B(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6742_ (.A1(_1971_),
    .A2(_2060_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6743_ (.A1(_1000_),
    .A2(_1908_),
    .B(_1810_),
    .C(_2061_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6744_ (.A1(_0553_),
    .A2(_1966_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6745_ (.A1(_1808_),
    .A2(_2062_),
    .A3(_2063_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6746_ (.A1(_0516_),
    .A2(_2056_),
    .B(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6747_ (.A1(_0511_),
    .A2(_1832_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6748_ (.A1(_1803_),
    .A2(_2065_),
    .B(_2066_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6749_ (.A1(_2013_),
    .A2(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6750_ (.I(_1864_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6751_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6752_ (.I(_1801_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6753_ (.A1(_2049_),
    .A2(_2052_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6754_ (.A1(_2034_),
    .A2(_2047_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6755_ (.A1(_1987_),
    .A2(_2048_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6756_ (.A1(_2073_),
    .A2(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6757_ (.I(_1936_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6758_ (.A1(_0517_),
    .A2(_2076_),
    .A3(_2045_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6759_ (.A1(_2040_),
    .A2(_2044_),
    .B(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6760_ (.A1(_2037_),
    .A2(_2042_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6761_ (.A1(_2041_),
    .A2(_2043_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6762_ (.A1(_2079_),
    .A2(_2080_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6763_ (.A1(_0710_),
    .A2(_2036_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6764_ (.A1(_4209_),
    .A2(_0526_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6765_ (.A1(_2082_),
    .A2(_2083_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6766_ (.A1(_2082_),
    .A2(_2083_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6767_ (.A1(_2084_),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6768_ (.A1(_2081_),
    .A2(_2086_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6769_ (.A1(_1937_),
    .A2(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6770_ (.A1(_2078_),
    .A2(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6771_ (.A1(_2075_),
    .A2(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6772_ (.A1(_2028_),
    .A2(_2053_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6773_ (.A1(_2028_),
    .A2(_2029_),
    .B(_2053_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6774_ (.A1(_2006_),
    .A2(_2009_),
    .A3(_2091_),
    .B(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6775_ (.A1(_2072_),
    .A2(_2090_),
    .A3(_2093_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6776_ (.A1(_2071_),
    .A2(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6777_ (.A1(_1962_),
    .A2(_2068_),
    .B(_2070_),
    .C(_2095_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6778_ (.I(_0649_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6779_ (.A1(_0607_),
    .A2(_1853_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6780_ (.A1(_1281_),
    .A2(_1910_),
    .B(_2097_),
    .C(_1836_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6781_ (.A1(_0602_),
    .A2(_1968_),
    .B(_1838_),
    .C(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6782_ (.A1(_0591_),
    .A2(_1909_),
    .B(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6783_ (.A1(_1971_),
    .A2(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6784_ (.A1(_1022_),
    .A2(_1908_),
    .B(_1829_),
    .C(_2101_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6785_ (.A1(_0587_),
    .A2(_1966_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6786_ (.A1(_1808_),
    .A2(_2102_),
    .A3(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6787_ (.A1(_0619_),
    .A2(_2056_),
    .B(_1832_),
    .C(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6788_ (.A1(_2096_),
    .A2(_1803_),
    .B(_2105_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6789_ (.A1(_1964_),
    .A2(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6790_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_2069_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6791_ (.A1(_2072_),
    .A2(_2090_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6792_ (.A1(_2072_),
    .A2(_2090_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6793_ (.A1(_2109_),
    .A2(_2093_),
    .B(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6794_ (.A1(_0588_),
    .A2(_2076_),
    .A3(_2087_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6795_ (.A1(_2081_),
    .A2(_2086_),
    .B(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6796_ (.A1(_0710_),
    .A2(_2076_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6797_ (.A1(_4210_),
    .A2(_2036_),
    .A3(_2042_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6798_ (.A1(_2114_),
    .A2(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6799_ (.I(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6800_ (.A1(_2113_),
    .A2(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6801_ (.I(_2078_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6802_ (.A1(_2119_),
    .A2(_2088_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6803_ (.A1(_2073_),
    .A2(_2074_),
    .B(_2089_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6804_ (.A1(_2120_),
    .A2(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6805_ (.A1(_2118_),
    .A2(_2122_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6806_ (.A1(_2111_),
    .A2(_2123_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6807_ (.A1(_2071_),
    .A2(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6808_ (.A1(_1962_),
    .A2(_2107_),
    .B(_2108_),
    .C(_2125_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6809_ (.A1(_2121_),
    .A2(_2118_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6810_ (.A1(_2111_),
    .A2(_2123_),
    .B(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6811_ (.A1(_1986_),
    .A2(_2082_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6812_ (.A1(_1986_),
    .A2(_2084_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6813_ (.A1(_2128_),
    .A2(_2129_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6814_ (.A1(_2113_),
    .A2(_2117_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6815_ (.A1(_2120_),
    .A2(_2118_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6816_ (.A1(_2131_),
    .A2(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6817_ (.A1(_2130_),
    .A2(_2133_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6818_ (.A1(_2127_),
    .A2(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6819_ (.A1(_0680_),
    .A2(_0720_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6820_ (.A1(_2136_),
    .A2(_1853_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6821_ (.A1(_1373_),
    .A2(_1823_),
    .B(_2137_),
    .C(_1836_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6822_ (.A1(_4223_),
    .A2(_1968_),
    .B(_1818_),
    .C(_2138_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6823_ (.A1(_0646_),
    .A2(_1819_),
    .B(_2139_),
    .C(_1815_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6824_ (.A1(_0712_),
    .A2(_1971_),
    .B(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6825_ (.A1(_1810_),
    .A2(_2141_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6826_ (.A1(_0709_),
    .A2(_1918_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6827_ (.A1(_1807_),
    .A2(_2142_),
    .A3(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6828_ (.A1(_0735_),
    .A2(_2056_),
    .B(_1848_),
    .C(_2144_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6829_ (.A1(_0701_),
    .A2(_1848_),
    .B(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6830_ (.A1(_1964_),
    .A2(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6831_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_2069_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6832_ (.A1(_2013_),
    .A2(_2135_),
    .B1(_2147_),
    .B2(_1852_),
    .C(_2148_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6833_ (.A1(_2127_),
    .A2(_2134_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6834_ (.A1(_2131_),
    .A2(_2132_),
    .B(_2129_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6835_ (.A1(_2128_),
    .A2(_2149_),
    .A3(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6836_ (.A1(_4225_),
    .A2(_0782_),
    .A3(_1813_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6837_ (.A1(_1519_),
    .A2(_1854_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6838_ (.A1(_0787_),
    .A2(_1855_),
    .B(_2153_),
    .C(_1821_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6839_ (.A1(_1819_),
    .A2(_2152_),
    .A3(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6840_ (.A1(_1386_),
    .A2(_1839_),
    .B(_2155_),
    .C(_1816_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6841_ (.A1(_1039_),
    .A2(_1908_),
    .B(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6842_ (.A1(_1844_),
    .A2(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6843_ (.A1(_0781_),
    .A2(_1810_),
    .B(_2056_),
    .C(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6844_ (.A1(_0797_),
    .A2(_1907_),
    .B(_1965_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6845_ (.A1(_0804_),
    .A2(_0815_),
    .B(_1832_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6846_ (.A1(_2159_),
    .A2(_2160_),
    .B(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6847_ (.A1(_1964_),
    .A2(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6848_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_2069_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6849_ (.A1(_2013_),
    .A2(_2151_),
    .B1(_2163_),
    .B2(_1852_),
    .C(_2164_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6850_ (.A1(_1051_),
    .A2(_1766_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6851_ (.I(_2165_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6852_ (.I(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6853_ (.A1(_1747_),
    .A2(_1298_),
    .A3(_1601_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6854_ (.I(_2168_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6855_ (.A1(_1713_),
    .A2(_0977_),
    .A3(_1750_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6856_ (.I(_2170_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6857_ (.A1(_1598_),
    .A2(_2169_),
    .B1(_2171_),
    .B2(\as2650.stack[0][0] ),
    .C(_2166_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6858_ (.A1(_1590_),
    .A2(_2167_),
    .B(_2172_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6859_ (.A1(_1670_),
    .A2(_2169_),
    .B1(_2171_),
    .B2(\as2650.stack[0][1] ),
    .C(_2166_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6860_ (.A1(_1611_),
    .A2(_2167_),
    .B(_2173_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6861_ (.I(_2165_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6862_ (.A1(_1624_),
    .A2(_2169_),
    .B1(_2171_),
    .B2(\as2650.stack[0][2] ),
    .C(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6863_ (.A1(_1620_),
    .A2(_2167_),
    .B(_2175_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6864_ (.A1(_1632_),
    .A2(_2169_),
    .B1(_2171_),
    .B2(\as2650.stack[0][3] ),
    .C(_2174_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6865_ (.A1(_1727_),
    .A2(_2167_),
    .B(_2176_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6866_ (.I(_1635_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6867_ (.I(_2166_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6868_ (.I(_2168_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6869_ (.I(_2170_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6870_ (.A1(_1639_),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\as2650.stack[0][4] ),
    .C(_2174_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6871_ (.A1(_2177_),
    .A2(_2178_),
    .B(_2181_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6872_ (.A1(_1646_),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\as2650.stack[0][5] ),
    .C(_2174_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6873_ (.A1(_1642_),
    .A2(_2178_),
    .B(_2182_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6874_ (.A1(_1651_),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\as2650.stack[0][6] ),
    .C(_2165_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6875_ (.A1(_1649_),
    .A2(_2178_),
    .B(_2183_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6876_ (.A1(_1741_),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\as2650.stack[0][7] ),
    .C(_2165_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6877_ (.A1(_1698_),
    .A2(_2178_),
    .B(_2184_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6878_ (.A1(_1542_),
    .A2(_1850_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6879_ (.I(_2185_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6880_ (.A1(_1542_),
    .A2(_1862_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6881_ (.A1(_1800_),
    .A2(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6882_ (.I(_2188_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6883_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6884_ (.A1(_4306_),
    .A2(_4322_),
    .A3(_2071_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6885_ (.A1(_1835_),
    .A2(_2186_),
    .B(_2190_),
    .C(_2191_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6886_ (.I(_2185_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6887_ (.I(_2188_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6888_ (.A1(_0287_),
    .A2(_1905_),
    .B1(_2193_),
    .B2(\as2650.r123_2[1][1] ),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6889_ (.A1(_1923_),
    .A2(_2192_),
    .B(_2194_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6890_ (.A1(\as2650.r123_2[1][2] ),
    .A2(_2193_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6891_ (.A1(_0380_),
    .A2(_2071_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6892_ (.A1(_1979_),
    .A2(_2186_),
    .B(_2195_),
    .C(_2196_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6893_ (.A1(_0483_),
    .A2(_2012_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6894_ (.A1(\as2650.r123_2[1][3] ),
    .A2(_2189_),
    .B(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6895_ (.A1(_2026_),
    .A2(_2192_),
    .B(_2198_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6896_ (.A1(_0577_),
    .A2(_2012_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6897_ (.A1(\as2650.r123_2[1][4] ),
    .A2(_2189_),
    .B(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6898_ (.A1(_2068_),
    .A2(_2192_),
    .B(_2200_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6899_ (.A1(_0677_),
    .A2(_1905_),
    .B1(_2193_),
    .B2(\as2650.r123_2[1][5] ),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6900_ (.A1(_2107_),
    .A2(_2192_),
    .B(_2201_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6901_ (.A1(_0774_),
    .A2(_1905_),
    .B1(_2193_),
    .B2(\as2650.r123_2[1][6] ),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6902_ (.A1(_2147_),
    .A2(_2186_),
    .B(_2202_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6903_ (.A1(_0857_),
    .A2(_2012_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6904_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_2189_),
    .B(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6905_ (.A1(_2163_),
    .A2(_2186_),
    .B(_2204_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6906_ (.A1(_1842_),
    .A2(_1911_),
    .A3(_1829_),
    .A4(_1802_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6907_ (.A1(_4086_),
    .A2(_1806_),
    .B(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6908_ (.A1(_0945_),
    .A2(_2206_),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6909_ (.I(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6910_ (.A1(_0939_),
    .A2(_1096_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6911_ (.I(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6912_ (.A1(\as2650.r123_2[0][0] ),
    .A2(_2208_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6913_ (.A1(_0888_),
    .A2(_1096_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6914_ (.I(_2212_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6915_ (.A1(_0876_),
    .A2(_1799_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6916_ (.A1(_0925_),
    .A2(_2212_),
    .B(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6917_ (.A1(_1589_),
    .A2(_2213_),
    .B(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6918_ (.A1(_2210_),
    .A2(_2211_),
    .B(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6919_ (.A1(_1834_),
    .A2(_2208_),
    .B(_2217_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6920_ (.A1(_0965_),
    .A2(_1799_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6921_ (.I(_2218_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6922_ (.A1(_1777_),
    .A2(_2219_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6923_ (.I(_2214_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6924_ (.A1(_0959_),
    .A2(_2213_),
    .B(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6925_ (.A1(_0945_),
    .A2(_1850_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6926_ (.I(_2223_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6927_ (.A1(_1922_),
    .A2(_2208_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6928_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_2224_),
    .B(_2225_),
    .C(_2210_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6929_ (.A1(_2220_),
    .A2(_2222_),
    .B(_2226_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6930_ (.I(_2209_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6931_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_2224_),
    .B(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6932_ (.I(_2207_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6933_ (.A1(_1978_),
    .A2(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6934_ (.I(_2218_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6935_ (.A1(_0980_),
    .A2(_2219_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6936_ (.A1(_0981_),
    .A2(_2231_),
    .B(_2221_),
    .C(_2232_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6937_ (.A1(_2228_),
    .A2(_2230_),
    .B(_2233_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6938_ (.A1(_0415_),
    .A2(_2219_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6939_ (.A1(_0994_),
    .A2(_2213_),
    .B(_2221_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6940_ (.A1(_2023_),
    .A2(_2024_),
    .A3(_2208_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6941_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_2224_),
    .B(_2236_),
    .C(_2210_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6942_ (.A1(_2234_),
    .A2(_2235_),
    .B(_2237_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6943_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_2224_),
    .B(_2227_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6944_ (.A1(_2067_),
    .A2(_2229_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6945_ (.A1(_1008_),
    .A2(_2218_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6946_ (.A1(_1000_),
    .A2(_2231_),
    .B(_2214_),
    .C(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6947_ (.A1(_2238_),
    .A2(_2239_),
    .B(_2241_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6948_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_2223_),
    .B(_2209_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6949_ (.A1(_2106_),
    .A2(_2229_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6950_ (.A1(_1021_),
    .A2(_2218_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6951_ (.A1(_1022_),
    .A2(_2231_),
    .B(_2214_),
    .C(_2244_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6952_ (.A1(_2242_),
    .A2(_2243_),
    .B(_2245_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6953_ (.A1(_1028_),
    .A2(_2219_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6954_ (.A1(_1034_),
    .A2(_2213_),
    .B(_2221_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6955_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_2223_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6956_ (.A1(_2146_),
    .A2(_2229_),
    .B(_2227_),
    .C(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6957_ (.A1(_2246_),
    .A2(_2247_),
    .B(_2249_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6958_ (.A1(\as2650.r123_2[0][7] ),
    .A2(_2223_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6959_ (.A1(_2162_),
    .A2(_2207_),
    .B(_2227_),
    .C(_2250_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6960_ (.A1(_1653_),
    .A2(_2231_),
    .A3(_2210_),
    .B(_2251_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6961_ (.I(\as2650.addr_buff[0] ),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6962_ (.A1(_1846_),
    .A2(_1543_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6963_ (.A1(_1445_),
    .A2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6964_ (.I(_4092_),
    .Z(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6965_ (.I(_2255_),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6966_ (.A1(_1241_),
    .A2(_1078_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6967_ (.A1(_1352_),
    .A2(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6968_ (.A1(_1258_),
    .A2(_2256_),
    .B1(_2258_),
    .B2(_1359_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6969_ (.I(_1072_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6970_ (.I(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6971_ (.A1(_2261_),
    .A2(_1548_),
    .B(_1567_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6972_ (.I(_1070_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6973_ (.A1(_4044_),
    .A2(_1052_),
    .A3(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6974_ (.I(_1079_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6975_ (.A1(_1443_),
    .A2(_4123_),
    .A3(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6976_ (.I(_1421_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6977_ (.I(_1450_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6978_ (.I(_4051_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6979_ (.I(_1059_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6980_ (.A1(_4119_),
    .A2(_4118_),
    .A3(_1246_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6981_ (.A1(_4046_),
    .A2(_2270_),
    .A3(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6982_ (.A1(_2269_),
    .A2(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6983_ (.A1(_2268_),
    .A2(_2273_),
    .B(_1449_),
    .C(_4284_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6984_ (.I(_4053_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6985_ (.A1(_2275_),
    .A2(_1253_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6986_ (.A1(_1057_),
    .A2(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6987_ (.A1(_2267_),
    .A2(_1062_),
    .B(_2274_),
    .C(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6988_ (.A1(_2262_),
    .A2(_2264_),
    .A3(_2266_),
    .A4(_2278_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6989_ (.I(_4293_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6990_ (.A1(_1074_),
    .A2(_1077_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6991_ (.I(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6992_ (.A1(_4035_),
    .A2(_1062_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6993_ (.A1(_1567_),
    .A2(_2282_),
    .A3(_1430_),
    .A4(_2283_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6994_ (.A1(_4105_),
    .A2(_1845_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6995_ (.A1(_4047_),
    .A2(_4051_),
    .A3(_2270_),
    .A4(_2271_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6996_ (.A1(_4091_),
    .A2(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6997_ (.A1(_4029_),
    .A2(_1054_),
    .A3(_2275_),
    .A4(_4102_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6998_ (.A1(_2288_),
    .A2(_2272_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6999_ (.A1(_2285_),
    .A2(_2287_),
    .A3(_2289_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7000_ (.A1(_1426_),
    .A2(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7001_ (.A1(_2280_),
    .A2(_1548_),
    .A3(_2284_),
    .B(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7002_ (.A1(_2254_),
    .A2(_2259_),
    .A3(_2279_),
    .A4(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7003_ (.I(_2293_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7004_ (.I0(_2252_),
    .I1(_1559_),
    .S(_2294_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7005_ (.I(_2295_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7006_ (.I(\as2650.addr_buff[1] ),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7007_ (.I0(_2296_),
    .I1(_1572_),
    .S(_2294_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7008_ (.I(_2297_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7009_ (.I(\as2650.addr_buff[2] ),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7010_ (.I(_1405_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7011_ (.I0(_2298_),
    .I1(_2299_),
    .S(_2294_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7012_ (.I(_2300_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7013_ (.I(\as2650.addr_buff[3] ),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7014_ (.I(_2293_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7015_ (.I(_1407_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7016_ (.I(_2293_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7017_ (.A1(_2303_),
    .A2(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7018_ (.A1(_2301_),
    .A2(_2302_),
    .B(_2305_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _7019_ (.I(\as2650.addr_buff[4] ),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7020_ (.I(_1410_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7021_ (.A1(_2307_),
    .A2(_2304_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7022_ (.A1(_2306_),
    .A2(_2302_),
    .B(_2308_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7023_ (.A1(_1283_),
    .A2(_2304_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7024_ (.A1(_4266_),
    .A2(_2302_),
    .B(_2309_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7025_ (.A1(_1584_),
    .A2(_2304_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7026_ (.A1(_4268_),
    .A2(_2302_),
    .B(_2310_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7027_ (.I(_4093_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7028_ (.I(_2311_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7029_ (.I0(_2312_),
    .I1(_1586_),
    .S(_2294_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7030_ (.I(_2313_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7031_ (.A1(_1272_),
    .A2(_1421_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7032_ (.A1(_1336_),
    .A2(_1223_),
    .B(_1363_),
    .C(_1226_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7033_ (.A1(_1271_),
    .A2(_1278_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7034_ (.A1(_2316_),
    .A2(_1462_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7035_ (.A1(_1344_),
    .A2(_1460_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7036_ (.I(_2318_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7037_ (.I(_1845_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7038_ (.A1(_1254_),
    .A2(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7039_ (.A1(_2319_),
    .A2(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7040_ (.A1(_4035_),
    .A2(_1562_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7041_ (.A1(_1442_),
    .A2(_2323_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7042_ (.I(_2283_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7043_ (.A1(_4195_),
    .A2(_1368_),
    .A3(_2325_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7044_ (.A1(_2322_),
    .A2(_2324_),
    .A3(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7045_ (.A1(_1062_),
    .A2(_1431_),
    .B(_2317_),
    .C(_2327_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7046_ (.A1(_2314_),
    .A2(_2315_),
    .B(_2328_),
    .C(_2254_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7047_ (.A1(_4089_),
    .A2(_2283_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7048_ (.I(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7049_ (.A1(_1474_),
    .A2(_1249_),
    .B(_2331_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7050_ (.A1(net24),
    .A2(_2329_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7051_ (.A1(_2329_),
    .A2(_2332_),
    .B(_2333_),
    .C(_1295_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7052_ (.I(_1251_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7053_ (.I(_1272_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7054_ (.I(_2335_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7055_ (.A1(_2334_),
    .A2(_2336_),
    .A3(_1286_),
    .A4(_1223_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7056_ (.I(_4284_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7057_ (.I(_2338_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7058_ (.A1(net22),
    .A2(_2337_),
    .B(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7059_ (.A1(_4166_),
    .A2(_2337_),
    .B(_2340_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7060_ (.I(_1057_),
    .Z(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7061_ (.A1(_2275_),
    .A2(_2341_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7062_ (.I(_2276_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7063_ (.I(_2343_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7064_ (.A1(_1450_),
    .A2(_2343_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7065_ (.A1(_1272_),
    .A2(_2345_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7066_ (.A1(_2316_),
    .A2(_2344_),
    .B1(_2322_),
    .B2(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7067_ (.A1(_1253_),
    .A2(_1226_),
    .A3(_2314_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7068_ (.A1(_1394_),
    .A2(_1449_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7069_ (.A1(_1226_),
    .A2(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7070_ (.A1(_2344_),
    .A2(_2348_),
    .A3(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7071_ (.A1(_1252_),
    .A2(_1544_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7072_ (.I(_1428_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7073_ (.I(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7074_ (.A1(_1069_),
    .A2(_2318_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7075_ (.A1(_2354_),
    .A2(_2355_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7076_ (.A1(_2347_),
    .A2(_2351_),
    .A3(_2352_),
    .A4(_2356_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7077_ (.A1(net23),
    .A2(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7078_ (.A1(_2342_),
    .A2(_2357_),
    .B(_2358_),
    .C(_1471_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7079_ (.A1(_0868_),
    .A2(_1520_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7080_ (.I(_2359_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7081_ (.I(_2360_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7082_ (.I(_2359_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7083_ (.A1(_0940_),
    .A2(_4315_),
    .A3(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7084_ (.I(_2363_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7085_ (.A1(_4317_),
    .A2(_1903_),
    .B1(_2364_),
    .B2(\as2650.r123[2][0] ),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7086_ (.A1(_4283_),
    .A2(_2361_),
    .B(_2365_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7087_ (.A1(_4317_),
    .A2(_1960_),
    .B1(_2364_),
    .B2(\as2650.r123[2][1] ),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7088_ (.A1(_4412_),
    .A2(_2361_),
    .B(_2366_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7089_ (.A1(_4317_),
    .A2(_2010_),
    .B1(_2364_),
    .B2(\as2650.r123[2][2] ),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7090_ (.A1(_0366_),
    .A2(_2361_),
    .B(_2367_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7091_ (.I(_2363_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7092_ (.A1(_0288_),
    .A2(_2054_),
    .B1(_2368_),
    .B2(\as2650.r123[2][3] ),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7093_ (.A1(_0461_),
    .A2(_2361_),
    .B(_2369_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7094_ (.A1(_0288_),
    .A2(_2094_),
    .B1(_2368_),
    .B2(\as2650.r123[2][4] ),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7095_ (.A1(_0558_),
    .A2(_2360_),
    .B(_2370_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7096_ (.A1(_0288_),
    .A2(_2124_),
    .B1(_2368_),
    .B2(\as2650.r123[2][5] ),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7097_ (.A1(_0651_),
    .A2(_2360_),
    .B(_2371_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7098_ (.A1(\as2650.r123[2][6] ),
    .A2(_2364_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7099_ (.A1(_0462_),
    .A2(_2135_),
    .B1(_2360_),
    .B2(_0738_),
    .C(_2372_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7100_ (.A1(_0817_),
    .A2(_2362_),
    .B1(_2368_),
    .B2(\as2650.r123[2][7] ),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7101_ (.A1(_0462_),
    .A2(_2151_),
    .B(_2373_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7102_ (.A1(_4005_),
    .A2(_1451_),
    .A3(_1217_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7103_ (.A1(_1343_),
    .A2(_1452_),
    .A3(_1453_),
    .B(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7104_ (.A1(_4049_),
    .A2(_1561_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7105_ (.I(_0934_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7106_ (.A1(_4307_),
    .A2(_1436_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7107_ (.A1(_1284_),
    .A2(_2377_),
    .B(_2378_),
    .C(_2356_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7108_ (.A1(_1232_),
    .A2(_0874_),
    .A3(_1235_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7109_ (.A1(_1341_),
    .A2(_4170_),
    .A3(_1235_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7110_ (.A1(_2380_),
    .A2(_2381_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7111_ (.A1(_2258_),
    .A2(_2382_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7112_ (.A1(_1859_),
    .A2(_2376_),
    .B(_2379_),
    .C(_2383_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7113_ (.A1(_2347_),
    .A2(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7114_ (.A1(_4088_),
    .A2(_4027_),
    .A3(_4400_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7115_ (.I(_4250_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7116_ (.A1(_2387_),
    .A2(_0357_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7117_ (.A1(_0436_),
    .A2(_0543_),
    .A3(_0607_),
    .A4(_2388_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7118_ (.A1(_2136_),
    .A2(_0787_),
    .A3(_2386_),
    .A4(_2389_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7119_ (.A1(_2258_),
    .A2(_2390_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7120_ (.A1(_2375_),
    .A2(_2385_),
    .A3(_2391_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7121_ (.A1(_4364_),
    .A2(_2290_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7122_ (.A1(_1342_),
    .A2(_2277_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7123_ (.A1(_4038_),
    .A2(_1543_),
    .A3(_2289_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7124_ (.A1(_1429_),
    .A2(_2394_),
    .A3(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7125_ (.A1(_2393_),
    .A2(_2396_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7126_ (.A1(_4108_),
    .A2(_1219_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7127_ (.A1(_1554_),
    .A2(_1546_),
    .B(_2397_),
    .C(_2398_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7128_ (.A1(_4301_),
    .A2(_4084_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7129_ (.A1(\as2650.halted ),
    .A2(_1465_),
    .A3(_1543_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7130_ (.A1(_2400_),
    .A2(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7131_ (.A1(_4090_),
    .A2(_2270_),
    .A3(_2271_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7132_ (.A1(_2269_),
    .A2(_2403_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7133_ (.A1(_2286_),
    .A2(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7134_ (.A1(_1426_),
    .A2(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7135_ (.A1(_2268_),
    .A2(_1334_),
    .A3(_2257_),
    .A4(_2343_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7136_ (.I(_2269_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7137_ (.A1(_2408_),
    .A2(_2272_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7138_ (.I(_2394_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7139_ (.A1(_0785_),
    .A2(_2409_),
    .A3(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7140_ (.A1(_2407_),
    .A2(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7141_ (.A1(_2312_),
    .A2(_4261_),
    .B(_2331_),
    .C(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7142_ (.A1(_0965_),
    .A2(_2406_),
    .A3(_2413_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7143_ (.I(_1056_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7144_ (.I(_2415_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7145_ (.A1(_1074_),
    .A2(_1070_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7146_ (.A1(_0527_),
    .A2(_1451_),
    .A3(_1216_),
    .B1(_2417_),
    .B2(_1253_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7147_ (.A1(_1444_),
    .A2(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7148_ (.A1(_4362_),
    .A2(_2416_),
    .B(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7149_ (.A1(_1451_),
    .A2(_1423_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7150_ (.A1(_4049_),
    .A2(_1270_),
    .A3(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7151_ (.A1(_2343_),
    .A2(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7152_ (.A1(_1050_),
    .A2(_2423_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7153_ (.A1(_2402_),
    .A2(_2414_),
    .A3(_2420_),
    .A4(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7154_ (.A1(_2392_),
    .A2(_2399_),
    .A3(_2425_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7155_ (.I(_0883_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7156_ (.I(_2427_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7157_ (.A1(net54),
    .A2(_2428_),
    .B(_1459_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7158_ (.I(_1242_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7159_ (.I(_2430_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7160_ (.A1(_4070_),
    .A2(_1348_),
    .B(_1460_),
    .C(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7161_ (.I(_2265_),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7162_ (.I(_2433_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7163_ (.A1(net54),
    .A2(_2428_),
    .A3(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7164_ (.A1(_2429_),
    .A2(_2432_),
    .B(_2435_),
    .C(_1362_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7165_ (.A1(_1358_),
    .A2(_2323_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7166_ (.I(_2437_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7167_ (.I(_4194_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7168_ (.I(_1063_),
    .Z(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7169_ (.A1(_2341_),
    .A2(_1552_),
    .B1(_2439_),
    .B2(net54),
    .C(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7170_ (.A1(_2438_),
    .A2(_2441_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7171_ (.A1(_2436_),
    .A2(_2442_),
    .B(_2426_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7172_ (.A1(net49),
    .A2(_2426_),
    .B(_2443_),
    .C(_1295_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7173_ (.A1(_1224_),
    .A2(_2353_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7174_ (.I(_2444_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7175_ (.I(_2445_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7176_ (.A1(_1251_),
    .A2(_0888_),
    .A3(_1094_),
    .A4(_1465_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7177_ (.A1(_1568_),
    .A2(_2446_),
    .B(_2447_),
    .C(_2418_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7178_ (.A1(_4036_),
    .A2(_4122_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7179_ (.A1(_2282_),
    .A2(_2449_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7180_ (.A1(_1271_),
    .A2(_4089_),
    .A3(_1552_),
    .A4(_4123_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7181_ (.A1(_2450_),
    .A2(_2451_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7182_ (.A1(_4054_),
    .A2(_4122_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7183_ (.A1(_4301_),
    .A2(_4084_),
    .B1(_1079_),
    .B2(_2453_),
    .C(_2398_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7184_ (.A1(_2392_),
    .A2(_2448_),
    .A3(_2452_),
    .A4(_2454_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7185_ (.A1(net25),
    .A2(_1553_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7186_ (.A1(_1064_),
    .A2(_2456_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7187_ (.A1(_2427_),
    .A2(_2410_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7188_ (.I(_2458_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7189_ (.A1(_1421_),
    .A2(_2277_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7190_ (.I(_2460_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7191_ (.I(_2461_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7192_ (.A1(_1459_),
    .A2(_1460_),
    .B(_2456_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7193_ (.I(_1546_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7194_ (.I(_2464_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7195_ (.I(_2282_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7196_ (.A1(_2260_),
    .A2(_2466_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7197_ (.A1(_1066_),
    .A2(_2465_),
    .A3(_2456_),
    .A4(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7198_ (.I(_2417_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7199_ (.I(_2469_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7200_ (.A1(_1242_),
    .A2(_4292_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7201_ (.I(_2471_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7202_ (.I(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7203_ (.A1(_1523_),
    .A2(_2470_),
    .B(_2473_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7204_ (.A1(_2336_),
    .A2(_1348_),
    .A3(_2463_),
    .B1(_2468_),
    .B2(_2474_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7205_ (.A1(_2462_),
    .A2(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7206_ (.A1(_2457_),
    .A2(_2459_),
    .B(_1563_),
    .C(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7207_ (.A1(net25),
    .A2(_2455_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7208_ (.I(_1294_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7209_ (.A1(_2455_),
    .A2(_2477_),
    .B(_2478_),
    .C(_2479_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7210_ (.I(_2345_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7211_ (.I(_2267_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7212_ (.I(_2255_),
    .Z(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7213_ (.A1(_2481_),
    .A2(_1552_),
    .A3(_2482_),
    .A4(_2325_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7214_ (.A1(_1445_),
    .A2(_2480_),
    .A3(_2395_),
    .A4(_2483_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7215_ (.I(_2323_),
    .Z(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7216_ (.A1(_4095_),
    .A2(_2485_),
    .B(_2484_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7217_ (.A1(_4058_),
    .A2(_2484_),
    .B(_2486_),
    .C(_2479_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7218_ (.A1(_4094_),
    .A2(_2485_),
    .B(_2484_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7219_ (.A1(_4057_),
    .A2(_2484_),
    .B(_2487_),
    .C(_2479_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7220_ (.A1(_4189_),
    .A2(_1317_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7221_ (.I(_0937_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7222_ (.I(_2489_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7223_ (.A1(_1399_),
    .A2(_2490_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7224_ (.A1(_2488_),
    .A2(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7225_ (.I(_0640_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7226_ (.I(_1462_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7227_ (.A1(_1214_),
    .A2(_0397_),
    .A3(_1345_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7228_ (.A1(_1358_),
    .A2(_1551_),
    .A3(_1562_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7229_ (.A1(_1797_),
    .A2(_1436_),
    .B(_1440_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7230_ (.A1(_4194_),
    .A2(_1454_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7231_ (.A1(_2495_),
    .A2(_2496_),
    .A3(_2497_),
    .A4(_2498_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7232_ (.A1(_2493_),
    .A2(_2494_),
    .B(_2499_),
    .C(_1465_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7233_ (.I(_2500_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7234_ (.I0(\as2650.holding_reg[0] ),
    .I1(_2492_),
    .S(_2501_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7235_ (.I(_2502_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7236_ (.I(_2500_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7237_ (.I(_2490_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7238_ (.A1(_1401_),
    .A2(_1355_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7239_ (.I(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7240_ (.A1(_1777_),
    .A2(_2504_),
    .B(_2506_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7241_ (.A1(_4326_),
    .A2(_2503_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7242_ (.A1(_2503_),
    .A2(_2507_),
    .B(_2508_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7243_ (.A1(_0981_),
    .A2(_1348_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7244_ (.A1(_2299_),
    .A2(_1286_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7245_ (.A1(_2509_),
    .A2(_2510_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7246_ (.I0(_0387_),
    .I1(_2511_),
    .S(_2501_),
    .Z(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7247_ (.I(_2512_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7248_ (.I(_2280_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7249_ (.A1(_1407_),
    .A2(_2513_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7250_ (.A1(_1627_),
    .A2(_2513_),
    .B(_2514_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7251_ (.I0(_0395_),
    .I1(_2515_),
    .S(_2501_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7252_ (.I(_2516_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7253_ (.I(_1481_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7254_ (.A1(_2307_),
    .A2(_2513_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7255_ (.A1(_1635_),
    .A2(_2517_),
    .B(_2518_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7256_ (.I0(_0490_),
    .I1(_2519_),
    .S(_2501_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7257_ (.I(_2520_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7258_ (.A1(_1282_),
    .A2(_2489_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7259_ (.A1(_1280_),
    .A2(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7260_ (.I0(_0636_),
    .I1(_2522_),
    .S(_2500_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7261_ (.I(_2523_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7262_ (.A1(_1028_),
    .A2(_1286_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7263_ (.A1(_1584_),
    .A2(_2513_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7264_ (.A1(_2524_),
    .A2(_2525_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7265_ (.I0(_0689_),
    .I1(_2526_),
    .S(_2500_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7266_ (.I(_2527_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7267_ (.A1(_1523_),
    .A2(_2517_),
    .B(_1526_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7268_ (.A1(_2503_),
    .A2(_2528_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7269_ (.A1(_0799_),
    .A2(_2503_),
    .B(_2529_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7270_ (.I(_4287_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7271_ (.I(_2530_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7272_ (.I(_1293_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7273_ (.I(_2532_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7274_ (.A1(_2531_),
    .A2(_2378_),
    .B(_2533_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7275_ (.I(_4285_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7276_ (.A1(_2334_),
    .A2(_2534_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7277_ (.I(_1546_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7278_ (.A1(_2430_),
    .A2(_2536_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7279_ (.A1(_2382_),
    .A2(_2390_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7280_ (.A1(_4292_),
    .A2(_2538_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7281_ (.A1(_2341_),
    .A2(_2321_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7282_ (.A1(_1550_),
    .A2(_4122_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7283_ (.I(_1065_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7284_ (.A1(_2434_),
    .A2(_2542_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7285_ (.A1(_2434_),
    .A2(_2539_),
    .A3(_2540_),
    .B1(_2541_),
    .B2(_2543_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7286_ (.I(_2415_),
    .Z(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7287_ (.I(_2545_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7288_ (.I(_2546_),
    .Z(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7289_ (.I(_4081_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7290_ (.A1(_2341_),
    .A2(_2548_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7291_ (.I(_4079_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7292_ (.A1(_1260_),
    .A2(_1263_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7293_ (.A1(_1560_),
    .A2(_2550_),
    .A3(_2551_),
    .A4(_1229_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7294_ (.A1(_2547_),
    .A2(_2319_),
    .B1(_2549_),
    .B2(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7295_ (.A1(_1237_),
    .A2(_2549_),
    .B(_1230_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7296_ (.A1(_2553_),
    .A2(_2554_),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7297_ (.A1(_2537_),
    .A2(_2544_),
    .B1(_2555_),
    .B2(_2431_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7298_ (.A1(_2480_),
    .A2(_2556_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7299_ (.I(_0785_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7300_ (.I(_2409_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7301_ (.A1(_2558_),
    .A2(_2439_),
    .B(_2559_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7302_ (.A1(_4090_),
    .A2(_4056_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7303_ (.A1(_2311_),
    .A2(_2561_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7304_ (.A1(_4194_),
    .A2(_4056_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7305_ (.A1(_2562_),
    .A2(_2563_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7306_ (.A1(_2326_),
    .A2(_2564_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7307_ (.A1(_4056_),
    .A2(_2540_),
    .B(_2560_),
    .C(_2565_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7308_ (.A1(_1578_),
    .A2(_1433_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7309_ (.A1(_2481_),
    .A2(_2344_),
    .A3(_2566_),
    .A4(_2567_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7310_ (.A1(_1560_),
    .A2(_2464_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7311_ (.A1(_2534_),
    .A2(_2352_),
    .A3(_2568_),
    .A4(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7312_ (.A1(_1550_),
    .A2(_2535_),
    .B1(_2557_),
    .B2(_2570_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7313_ (.I(_2277_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7314_ (.I(_2571_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7315_ (.A1(_2263_),
    .A2(_2539_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7316_ (.A1(_4036_),
    .A2(_4054_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7317_ (.A1(_1549_),
    .A2(_2450_),
    .B(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7318_ (.I(_2466_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7319_ (.A1(_1257_),
    .A2(_2576_),
    .A3(_2440_),
    .A4(_2574_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7320_ (.A1(_2573_),
    .A2(_2575_),
    .A3(_2577_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7321_ (.I(_2574_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7322_ (.I(_2273_),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7323_ (.A1(_2579_),
    .A2(_2564_),
    .B(_2580_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7324_ (.A1(_2428_),
    .A2(_2440_),
    .A3(_2560_),
    .A4(_2581_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7325_ (.A1(_2344_),
    .A2(_2567_),
    .A3(_2582_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7326_ (.A1(_1230_),
    .A2(_1237_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7327_ (.A1(_1257_),
    .A2(_2574_),
    .B1(_2552_),
    .B2(_1481_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7328_ (.I(_1449_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7329_ (.A1(_2584_),
    .A2(_2585_),
    .B(_2586_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7330_ (.A1(_1569_),
    .A2(_2578_),
    .B1(_2583_),
    .B2(_2480_),
    .C(_2587_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7331_ (.A1(_1551_),
    .A2(_2572_),
    .A3(_2588_),
    .B1(_2535_),
    .B2(_2275_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7332_ (.I(_1252_),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7333_ (.I(_1293_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7334_ (.I(_2461_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7335_ (.I(_2464_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7336_ (.I(_2320_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7337_ (.I(_2593_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7338_ (.A1(_4121_),
    .A2(_4103_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7339_ (.A1(_2594_),
    .A2(_2595_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7340_ (.A1(_2449_),
    .A2(_2596_),
    .B(_2434_),
    .C(_2542_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7341_ (.A1(_1577_),
    .A2(_2353_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7342_ (.I(_2598_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7343_ (.I(_2466_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7344_ (.A1(_1249_),
    .A2(_2596_),
    .B(_2599_),
    .C(_2600_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7345_ (.A1(_1055_),
    .A2(_2592_),
    .B1(_2597_),
    .B2(_2601_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7346_ (.I(_1273_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7347_ (.A1(_1438_),
    .A2(_1230_),
    .B(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7348_ (.A1(_1430_),
    .A2(_2319_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7349_ (.I(_1439_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7350_ (.A1(_2550_),
    .A2(_2606_),
    .B(_2595_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7351_ (.A1(_2605_),
    .A2(_2607_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7352_ (.A1(_2336_),
    .A2(_2602_),
    .B1(_2604_),
    .B2(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7353_ (.A1(_2439_),
    .A2(_1346_),
    .A3(_1452_),
    .B(_2596_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7354_ (.I(_2410_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7355_ (.A1(_2591_),
    .A2(_2609_),
    .B1(_2610_),
    .B2(_2611_),
    .C(_2334_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7356_ (.A1(_2589_),
    .A2(_1054_),
    .B(_2590_),
    .C(_2612_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7357_ (.A1(_4029_),
    .A2(_4121_),
    .A3(_4103_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7358_ (.A1(_1054_),
    .A2(_1247_),
    .B(_1058_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7359_ (.A1(_2613_),
    .A2(_2614_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7360_ (.A1(_1064_),
    .A2(_2257_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7361_ (.A1(_2615_),
    .A2(_2616_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7362_ (.A1(_0784_),
    .A2(_2353_),
    .A3(_1545_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7363_ (.A1(_2542_),
    .A2(_1071_),
    .B(_2617_),
    .C(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7364_ (.I(_2559_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7365_ (.A1(_2439_),
    .A2(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7366_ (.I(_2255_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7367_ (.I(_2622_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7368_ (.A1(_2623_),
    .A2(_2563_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7369_ (.I(_2561_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7370_ (.I(_2625_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7371_ (.A1(_1231_),
    .A2(_2312_),
    .A3(_4074_),
    .B(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7372_ (.A1(_2624_),
    .A2(_2615_),
    .B(_2627_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7373_ (.I(_2273_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7374_ (.A1(_1523_),
    .A2(_2629_),
    .B(_2410_),
    .C(_2440_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7375_ (.A1(_2621_),
    .A2(_2628_),
    .B(_2630_),
    .C(_2326_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7376_ (.A1(_2591_),
    .A2(_2619_),
    .B(_2631_),
    .C(_2589_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7377_ (.A1(_2589_),
    .A2(_1058_),
    .B(_2590_),
    .C(_2632_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7378_ (.I(\as2650.cycle[4] ),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7379_ (.A1(_1252_),
    .A2(_2613_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7380_ (.A1(_2633_),
    .A2(_2634_),
    .B(_2339_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7381_ (.A1(_2633_),
    .A2(_2634_),
    .B(_2635_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7382_ (.A1(_4050_),
    .A2(_2633_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7383_ (.A1(_2613_),
    .A2(_2636_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7384_ (.A1(_2633_),
    .A2(_2634_),
    .B(_4050_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7385_ (.A1(_2531_),
    .A2(_2637_),
    .B(_2638_),
    .C(_2479_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7386_ (.I(_1293_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7387_ (.I(_2639_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7388_ (.A1(_2408_),
    .A2(_2637_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7389_ (.A1(_2408_),
    .A2(_2637_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7390_ (.A1(_4364_),
    .A2(_2580_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7391_ (.A1(_1843_),
    .A2(_2643_),
    .B(_2611_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7392_ (.A1(_2641_),
    .A2(_2642_),
    .A3(_2644_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7393_ (.A1(_2430_),
    .A2(_1334_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7394_ (.I(_2646_),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7395_ (.A1(_1578_),
    .A2(_2647_),
    .A3(_2611_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7396_ (.A1(_2531_),
    .A2(_2411_),
    .A3(_2645_),
    .A4(_2648_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7397_ (.A1(_2531_),
    .A2(_2408_),
    .B(_2649_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7398_ (.A1(_2640_),
    .A2(_2650_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7399_ (.I(_2494_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7400_ (.A1(_4128_),
    .A2(_2273_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7401_ (.A1(_4261_),
    .A2(_2651_),
    .A3(_2652_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7402_ (.A1(_4048_),
    .A2(_2641_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7403_ (.A1(_2647_),
    .A2(_2611_),
    .B1(_2653_),
    .B2(_2654_),
    .C(_2334_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7404_ (.A1(_2589_),
    .A2(_4048_),
    .B(_2590_),
    .C(_2655_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7405_ (.I(_4131_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7406_ (.A1(_2656_),
    .A2(_1370_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7407_ (.A1(_1500_),
    .A2(_2354_),
    .A3(_1370_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7408_ (.A1(_1487_),
    .A2(_1586_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7409_ (.A1(_1586_),
    .A2(_2657_),
    .B(_2658_),
    .C(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7410_ (.A1(_2374_),
    .A2(_2658_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7411_ (.A1(_1039_),
    .A2(_2374_),
    .B1(_2661_),
    .B2(net4),
    .C(_0861_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7412_ (.A1(_1487_),
    .A2(_2535_),
    .B1(_2660_),
    .B2(_2662_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7413_ (.A1(_2375_),
    .A2(_2420_),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7414_ (.A1(_1858_),
    .A2(_2355_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7415_ (.A1(_1463_),
    .A2(_2276_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7416_ (.A1(_2345_),
    .A2(_2664_),
    .B(_2665_),
    .C(_0876_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7417_ (.A1(_1240_),
    .A2(_1433_),
    .A3(_2380_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7418_ (.A1(_1417_),
    .A2(_4081_),
    .A3(_1545_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7419_ (.A1(_1845_),
    .A2(_2281_),
    .A3(_2288_),
    .A4(_2668_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7420_ (.A1(_2376_),
    .A2(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7421_ (.A1(_2396_),
    .A2(_2454_),
    .A3(_2667_),
    .A4(_2670_),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7422_ (.A1(_1065_),
    .A2(_2325_),
    .B(_1071_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7423_ (.A1(_1342_),
    .A2(_1063_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7424_ (.A1(_4362_),
    .A2(_2672_),
    .B(_2673_),
    .C(_2652_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7425_ (.A1(_1417_),
    .A2(_1229_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7426_ (.I(_2675_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7427_ (.A1(_1450_),
    .A2(_1091_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7428_ (.A1(_2676_),
    .A2(_2677_),
    .A3(_1561_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7429_ (.A1(_1437_),
    .A2(_2331_),
    .A3(_2678_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7430_ (.A1(_2311_),
    .A2(_0290_),
    .A3(_2265_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7431_ (.A1(_2401_),
    .A2(_2452_),
    .A3(_2618_),
    .A4(_2680_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7432_ (.A1(_2671_),
    .A2(_2674_),
    .A3(_2679_),
    .A4(_2681_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7433_ (.A1(_2424_),
    .A2(_2663_),
    .A3(_2666_),
    .A4(_2682_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7434_ (.I(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7435_ (.I(_2684_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7436_ (.I(_2685_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7437_ (.I(_2437_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7438_ (.I(_2687_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7439_ (.I(_1423_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7440_ (.I(_2316_),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7441_ (.I(_1045_),
    .Z(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7442_ (.I(_2691_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7443_ (.A1(\as2650.stack[7][0] ),
    .A2(_1298_),
    .B1(_2692_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7444_ (.I(_1175_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7445_ (.I(_2694_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7446_ (.A1(\as2650.stack[4][0] ),
    .A2(_1194_),
    .B1(_2695_),
    .B2(\as2650.stack[5][0] ),
    .C(_0915_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7447_ (.I(_1297_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7448_ (.A1(\as2650.stack[3][0] ),
    .A2(_2697_),
    .B1(_2692_),
    .B2(\as2650.stack[2][0] ),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7449_ (.A1(\as2650.stack[0][0] ),
    .A2(_1194_),
    .B1(_2695_),
    .B2(\as2650.stack[1][0] ),
    .C(_0923_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7450_ (.A1(_2693_),
    .A2(_2696_),
    .B1(_2698_),
    .B2(_2699_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7451_ (.I(_2469_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7452_ (.A1(_1597_),
    .A2(_1577_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7453_ (.A1(_1596_),
    .A2(_4062_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7454_ (.A1(_0937_),
    .A2(_2265_),
    .A3(_2538_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7455_ (.A1(_2702_),
    .A2(_2703_),
    .A3(_2704_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7456_ (.A1(_1254_),
    .A2(_2282_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7457_ (.A1(_2539_),
    .A2(_2706_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7458_ (.I(_1079_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7459_ (.A1(_4243_),
    .A2(_2415_),
    .B1(_2285_),
    .B2(\as2650.addr_buff[0] ),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7460_ (.A1(_1240_),
    .A2(_1443_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7461_ (.A1(\as2650.pc[0] ),
    .A2(net5),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7462_ (.A1(_1596_),
    .A2(_4242_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7463_ (.A1(_2711_),
    .A2(_2712_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7464_ (.A1(_2710_),
    .A2(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7465_ (.A1(_1597_),
    .A2(_2445_),
    .B(_2709_),
    .C(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7466_ (.A1(_4125_),
    .A2(_4151_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7467_ (.A1(_4242_),
    .A2(_2716_),
    .Z(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7468_ (.A1(_1439_),
    .A2(_2708_),
    .A3(_2717_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7469_ (.A1(_2708_),
    .A2(_2715_),
    .B(_2718_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7470_ (.A1(_1598_),
    .A2(_2707_),
    .B1(_2719_),
    .B2(_1797_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7471_ (.A1(_2705_),
    .A2(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7472_ (.A1(_2427_),
    .A2(_2713_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7473_ (.A1(_1666_),
    .A2(_1354_),
    .B(_2469_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7474_ (.I(_2430_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7475_ (.A1(_2701_),
    .A2(_2721_),
    .B1(_2722_),
    .B2(_2723_),
    .C(_2724_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7476_ (.A1(_1667_),
    .A2(_2689_),
    .B1(_2690_),
    .B2(_2700_),
    .C(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7477_ (.I(_2683_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7478_ (.A1(_2438_),
    .A2(_2726_),
    .B(_2727_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7479_ (.A1(_1765_),
    .A2(_2688_),
    .B(_2728_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7480_ (.I(_1294_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7481_ (.A1(_1765_),
    .A2(_2686_),
    .B(_2729_),
    .C(_2730_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7482_ (.I(_2727_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7483_ (.I(_2461_),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7484_ (.A1(_1612_),
    .A2(_1666_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7485_ (.I(_2733_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7486_ (.I(_1078_),
    .Z(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7487_ (.I(_2538_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7488_ (.A1(_2735_),
    .A2(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7489_ (.A1(_1613_),
    .A2(_2703_),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7490_ (.A1(_1481_),
    .A2(_2737_),
    .A3(_2738_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7491_ (.A1(_4241_),
    .A2(_4151_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7492_ (.A1(_1502_),
    .A2(_4233_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7493_ (.A1(_2740_),
    .A2(_2741_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7494_ (.A1(_1400_),
    .A2(_2416_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7495_ (.A1(_2594_),
    .A2(_2742_),
    .B(_2743_),
    .C(_2606_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7496_ (.A1(_1255_),
    .A2(_2708_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7497_ (.A1(_1550_),
    .A2(_2600_),
    .A3(_2734_),
    .B(_2745_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7498_ (.A1(_1335_),
    .A2(_2737_),
    .A3(_2734_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7499_ (.A1(\as2650.pc[1] ),
    .A2(net6),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7500_ (.A1(_2711_),
    .A2(_2748_),
    .Z(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7501_ (.A1(_4393_),
    .A2(_1072_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7502_ (.A1(\as2650.addr_buff[1] ),
    .A2(_2415_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7503_ (.A1(_1439_),
    .A2(_2750_),
    .A3(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7504_ (.A1(_2710_),
    .A2(_2749_),
    .B(_2752_),
    .C(_2263_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7505_ (.A1(_2445_),
    .A2(_2733_),
    .B(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7506_ (.A1(_2536_),
    .A2(_2749_),
    .B(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7507_ (.A1(_1354_),
    .A2(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7508_ (.A1(_2744_),
    .A2(_2746_),
    .B(_2747_),
    .C(_2756_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7509_ (.I(_2724_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7510_ (.A1(_2739_),
    .A2(_2757_),
    .B(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7511_ (.A1(_2724_),
    .A2(_1278_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7512_ (.A1(\as2650.stack[4][1] ),
    .A2(_1193_),
    .B1(_2694_),
    .B2(\as2650.stack[5][1] ),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7513_ (.I(_0911_),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7514_ (.A1(\as2650.stack[7][1] ),
    .A2(_2762_),
    .B1(_1046_),
    .B2(\as2650.stack[6][1] ),
    .C(_0913_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7515_ (.A1(\as2650.stack[3][1] ),
    .A2(_1296_),
    .B1(_1191_),
    .B2(\as2650.stack[0][1] ),
    .C1(\as2650.stack[1][1] ),
    .C2(_1175_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7516_ (.I(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7517_ (.A1(\as2650.stack[2][1] ),
    .A2(_2691_),
    .B(_2765_),
    .C(_0922_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7518_ (.A1(_2761_),
    .A2(_2763_),
    .B(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7519_ (.A1(_2316_),
    .A2(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7520_ (.A1(_2760_),
    .A2(_2734_),
    .B(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7521_ (.I(_2460_),
    .Z(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7522_ (.A1(_2759_),
    .A2(_2769_),
    .B(_2770_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7523_ (.A1(_2732_),
    .A2(_2734_),
    .B(_2771_),
    .C(_2727_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7524_ (.A1(_1615_),
    .A2(_2731_),
    .B(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7525_ (.A1(_2640_),
    .A2(_2773_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7526_ (.A1(_1679_),
    .A2(_2731_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7527_ (.I(_2684_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7528_ (.A1(_1612_),
    .A2(_1597_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7529_ (.A1(_1622_),
    .A2(_2776_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7530_ (.A1(_2539_),
    .A2(_2706_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7531_ (.I(_2778_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7532_ (.I(_2779_),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7533_ (.A1(_1353_),
    .A2(_1547_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7534_ (.I(_2781_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7535_ (.A1(\as2650.pc[1] ),
    .A2(net6),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7536_ (.A1(_2711_),
    .A2(_2748_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7537_ (.A1(_2783_),
    .A2(_2784_),
    .Z(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7538_ (.A1(\as2650.pc[2] ),
    .A2(_0347_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7539_ (.A1(_2785_),
    .A2(_2786_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7540_ (.A1(_1284_),
    .A2(_2536_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7541_ (.I(_1273_),
    .Z(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7542_ (.A1(_2782_),
    .A2(_2777_),
    .B1(_2787_),
    .B2(_2788_),
    .C(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7543_ (.I(_2460_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7544_ (.A1(_2780_),
    .A2(_2790_),
    .B(_2791_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7545_ (.A1(_0883_),
    .A2(_2736_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7546_ (.A1(_1613_),
    .A2(_2703_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7547_ (.A1(_1622_),
    .A2(_2794_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7548_ (.I(_2444_),
    .Z(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7549_ (.A1(_2796_),
    .A2(_2777_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7550_ (.A1(_2298_),
    .A2(_2545_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7551_ (.A1(_1575_),
    .A2(_2593_),
    .B(_1440_),
    .C(_2798_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7552_ (.A1(_1052_),
    .A2(_2787_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7553_ (.A1(_2797_),
    .A2(_2799_),
    .A3(_2800_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7554_ (.A1(_2793_),
    .A2(_2795_),
    .B1(_2801_),
    .B2(_2427_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7555_ (.I(_0290_),
    .Z(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7556_ (.I(_2803_),
    .Z(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7557_ (.A1(net7),
    .A2(_4384_),
    .Z(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7558_ (.A1(_4391_),
    .A2(_4233_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7559_ (.A1(_2740_),
    .A2(_2741_),
    .B(_2806_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7560_ (.A1(_2805_),
    .A2(_2807_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7561_ (.I(_2320_),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7562_ (.A1(_2805_),
    .A2(_2807_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7563_ (.A1(_2809_),
    .A2(_2810_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7564_ (.A1(_1575_),
    .A2(_2804_),
    .B1(_2808_),
    .B2(_2811_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7565_ (.I(_2745_),
    .Z(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7566_ (.A1(_2735_),
    .A2(_2802_),
    .B1(_2812_),
    .B2(_2813_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7567_ (.A1(_2592_),
    .A2(_2814_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7568_ (.A1(\as2650.stack[2][2] ),
    .A2(_2691_),
    .B1(_1193_),
    .B2(\as2650.stack[0][2] ),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7569_ (.A1(\as2650.stack[3][2] ),
    .A2(_1297_),
    .B1(_1176_),
    .B2(\as2650.stack[1][2] ),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7570_ (.A1(\as2650.stack[7][2] ),
    .A2(_2762_),
    .B1(_1046_),
    .B2(\as2650.stack[6][2] ),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7571_ (.I(_1191_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7572_ (.A1(\as2650.stack[4][2] ),
    .A2(_2819_),
    .B1(_2694_),
    .B2(\as2650.stack[5][2] ),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7573_ (.A1(_0922_),
    .A2(_2818_),
    .A3(_2820_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7574_ (.A1(_0914_),
    .A2(_2816_),
    .A3(_2817_),
    .B(_2821_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7575_ (.I(_2676_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7576_ (.I(_1423_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7577_ (.A1(_2824_),
    .A2(_2777_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7578_ (.A1(_2790_),
    .A2(_2815_),
    .B1(_2822_),
    .B2(_2823_),
    .C(_2825_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7579_ (.A1(_2777_),
    .A2(_2792_),
    .B1(_2826_),
    .B2(_2732_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7580_ (.A1(_2775_),
    .A2(_2827_),
    .B(_1471_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7581_ (.A1(_2774_),
    .A2(_2828_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7582_ (.I(_2683_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7583_ (.I(_2829_),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7584_ (.I(_2438_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7585_ (.I(_2824_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7586_ (.A1(\as2650.pc[2] ),
    .A2(\as2650.pc[1] ),
    .A3(\as2650.pc[0] ),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7587_ (.A1(_1630_),
    .A2(_2833_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7588_ (.A1(\as2650.stack[3][3] ),
    .A2(_2697_),
    .B1(_1047_),
    .B2(\as2650.stack[2][3] ),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7589_ (.I(_2819_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7590_ (.A1(\as2650.stack[0][3] ),
    .A2(_2836_),
    .B1(_2695_),
    .B2(\as2650.stack[1][3] ),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7591_ (.A1(\as2650.stack[7][3] ),
    .A2(_2697_),
    .B1(_1047_),
    .B2(\as2650.stack[6][3] ),
    .C1(_2836_),
    .C2(\as2650.stack[4][3] ),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7592_ (.A1(\as2650.stack[5][3] ),
    .A2(_1177_),
    .B(_0914_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7593_ (.A1(_0915_),
    .A2(_2835_),
    .A3(_2837_),
    .B1(_2838_),
    .B2(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7594_ (.I(_2840_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7595_ (.I(_2690_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7596_ (.I(_1052_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7597_ (.A1(_1630_),
    .A2(_0429_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7598_ (.A1(_1630_),
    .A2(net8),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7599_ (.A1(_2844_),
    .A2(_2845_),
    .Z(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7600_ (.A1(_1621_),
    .A2(_1402_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7601_ (.A1(_2785_),
    .A2(_2786_),
    .B(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7602_ (.A1(_2846_),
    .A2(_2848_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7603_ (.A1(_2843_),
    .A2(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7604_ (.I(_2260_),
    .Z(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7605_ (.A1(_1406_),
    .A2(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7606_ (.A1(_2301_),
    .A2(_2261_),
    .B(_2606_),
    .C(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7607_ (.A1(_2446_),
    .A2(_2834_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7608_ (.A1(_2850_),
    .A2(_2853_),
    .A3(_2854_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7609_ (.A1(_1336_),
    .A2(_2576_),
    .A3(_2855_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7610_ (.I(_2704_),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7611_ (.A1(_1621_),
    .A2(_1612_),
    .A3(_2703_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7612_ (.A1(_1631_),
    .A2(_2858_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7613_ (.I(_1072_),
    .Z(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7614_ (.I(_2860_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7615_ (.I(_2861_),
    .Z(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7616_ (.A1(_1402_),
    .A2(_4384_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7617_ (.A1(_0429_),
    .A2(_0340_),
    .Z(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7618_ (.A1(_2863_),
    .A2(_2810_),
    .B(_2864_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7619_ (.A1(_2863_),
    .A2(_2810_),
    .A3(_2864_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7620_ (.A1(_2862_),
    .A2(_2865_),
    .A3(_2866_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7621_ (.I(_2809_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7622_ (.I(_2745_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7623_ (.A1(_1406_),
    .A2(_2868_),
    .B(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7624_ (.A1(_2857_),
    .A2(_2859_),
    .B1(_2867_),
    .B2(_2870_),
    .C(_2465_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7625_ (.A1(_2647_),
    .A2(_2834_),
    .B1(_2849_),
    .B2(_2472_),
    .C(_2537_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7626_ (.A1(_2856_),
    .A2(_2871_),
    .B(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7627_ (.A1(_2832_),
    .A2(_2834_),
    .B1(_2841_),
    .B2(_2842_),
    .C(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7628_ (.A1(_2780_),
    .A2(_2872_),
    .B(_2791_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7629_ (.A1(_2834_),
    .A2(_2875_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7630_ (.A1(_2831_),
    .A2(_2874_),
    .B(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7631_ (.I(_2683_),
    .Z(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7632_ (.A1(_1729_),
    .A2(_2878_),
    .B(_2339_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7633_ (.A1(_2830_),
    .A2(_2877_),
    .B(_2879_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7634_ (.A1(_1684_),
    .A2(_2833_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7635_ (.A1(_1638_),
    .A2(_2880_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7636_ (.I(_2707_),
    .Z(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7637_ (.I(_2417_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7638_ (.I(_2883_),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7639_ (.A1(_1285_),
    .A2(_2884_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7640_ (.A1(_1687_),
    .A2(net9),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7641_ (.I(_2886_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7642_ (.I(_2845_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7643_ (.A1(_2844_),
    .A2(_2848_),
    .B(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7644_ (.A1(_2887_),
    .A2(_2889_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7645_ (.A1(_4307_),
    .A2(_2883_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7646_ (.I(_2891_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7647_ (.A1(_2885_),
    .A2(_2881_),
    .B1(_2890_),
    .B2(_2892_),
    .C(_2758_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7648_ (.I(_2687_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7649_ (.A1(_2882_),
    .A2(_2893_),
    .B(_2894_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7650_ (.A1(_1688_),
    .A2(_2880_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7651_ (.I(_2545_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7652_ (.I(_2897_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7653_ (.I(_0429_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7654_ (.A1(_2899_),
    .A2(_0340_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7655_ (.A1(net9),
    .A2(_0420_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7656_ (.I(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7657_ (.A1(_2900_),
    .A2(_2865_),
    .A3(_2902_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7658_ (.A1(_2900_),
    .A2(_2865_),
    .B(_2902_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7659_ (.A1(_1410_),
    .A2(_2593_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7660_ (.A1(_2898_),
    .A2(_2903_),
    .A3(_2904_),
    .B(_2905_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7661_ (.A1(_1683_),
    .A2(_2858_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7662_ (.A1(_1688_),
    .A2(_2907_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7663_ (.A1(_2793_),
    .A2(_2908_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7664_ (.A1(_1410_),
    .A2(_2809_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7665_ (.A1(\as2650.addr_buff[4] ),
    .A2(_2285_),
    .B1(_2598_),
    .B2(_2881_),
    .C1(_2890_),
    .C2(_2710_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7666_ (.A1(_2910_),
    .A2(_2911_),
    .B(_1335_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7667_ (.A1(_2909_),
    .A2(_2912_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7668_ (.A1(_2263_),
    .A2(_2913_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7669_ (.A1(_2813_),
    .A2(_2906_),
    .B(_2914_),
    .C(_2470_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7670_ (.A1(\as2650.stack[7][4] ),
    .A2(_2697_),
    .B1(_2836_),
    .B2(\as2650.stack[4][4] ),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7671_ (.A1(\as2650.stack[6][4] ),
    .A2(_2692_),
    .B1(_2695_),
    .B2(\as2650.stack[5][4] ),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7672_ (.A1(\as2650.stack[3][4] ),
    .A2(_1663_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7673_ (.A1(_0949_),
    .A2(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7674_ (.A1(\as2650.stack[0][4] ),
    .A2(_1193_),
    .B1(_1176_),
    .B2(\as2650.stack[1][4] ),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7675_ (.I(_2920_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7676_ (.A1(\as2650.stack[2][4] ),
    .A2(_2692_),
    .B(_2919_),
    .C(_2921_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7677_ (.A1(_0923_),
    .A2(_2916_),
    .A3(_2917_),
    .B(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7678_ (.A1(_2823_),
    .A2(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7679_ (.A1(_2689_),
    .A2(_2896_),
    .B1(_2893_),
    .B2(_2915_),
    .C(_2924_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7680_ (.A1(_2881_),
    .A2(_2895_),
    .B1(_2925_),
    .B2(_2688_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7681_ (.I(_2338_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7682_ (.A1(_1640_),
    .A2(_2878_),
    .B(_2927_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7683_ (.A1(_2830_),
    .A2(_2926_),
    .B(_2928_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7684_ (.A1(_1693_),
    .A2(_2878_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7685_ (.A1(_1688_),
    .A2(_1683_),
    .A3(_2833_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7686_ (.A1(_1643_),
    .A2(_2930_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _7687_ (.A1(\as2650.pc[5] ),
    .A2(net1),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7688_ (.A1(\as2650.pc[4] ),
    .A2(net9),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7689_ (.A1(_2887_),
    .A2(_2889_),
    .B(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7690_ (.A1(_2932_),
    .A2(_2934_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7691_ (.A1(_2891_),
    .A2(_2935_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7692_ (.A1(_2782_),
    .A2(_2931_),
    .B(_2936_),
    .C(_2603_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7693_ (.A1(_1638_),
    .A2(_2907_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7694_ (.A1(_1644_),
    .A2(_2938_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7695_ (.A1(_0538_),
    .A2(_0420_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7696_ (.A1(_0603_),
    .A2(_0531_),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7697_ (.A1(_2940_),
    .A2(_2904_),
    .A3(_2941_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7698_ (.A1(_2940_),
    .A2(_2904_),
    .B(_2941_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7699_ (.A1(_2851_),
    .A2(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7700_ (.A1(_2942_),
    .A2(_2944_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7701_ (.A1(_1287_),
    .A2(_2868_),
    .B(_2869_),
    .C(_2945_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7702_ (.I(_2710_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7703_ (.A1(_4095_),
    .A2(_2416_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7704_ (.A1(_1281_),
    .A2(_2860_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7705_ (.A1(_1440_),
    .A2(_2948_),
    .A3(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7706_ (.A1(_2947_),
    .A2(_2935_),
    .B(_2950_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7707_ (.A1(_2446_),
    .A2(_2931_),
    .B(_2951_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7708_ (.A1(_1317_),
    .A2(_2433_),
    .A3(_2952_),
    .B(_2884_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7709_ (.A1(_2857_),
    .A2(_2939_),
    .B(_2946_),
    .C(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7710_ (.A1(\as2650.stack[3][5] ),
    .A2(_2762_),
    .B1(_1045_),
    .B2(\as2650.stack[2][5] ),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7711_ (.I(_1175_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7712_ (.A1(\as2650.stack[0][5] ),
    .A2(_1192_),
    .B1(_2956_),
    .B2(\as2650.stack[1][5] ),
    .C(_0921_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7713_ (.A1(\as2650.stack[4][5] ),
    .A2(_1192_),
    .B1(_2956_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7714_ (.A1(\as2650.stack[7][5] ),
    .A2(_1296_),
    .B1(_1045_),
    .B2(\as2650.stack[6][5] ),
    .C(_0913_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7715_ (.A1(_2955_),
    .A2(_2957_),
    .B1(_2958_),
    .B2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7716_ (.I(_2823_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7717_ (.A1(_2824_),
    .A2(_2931_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7718_ (.A1(_2937_),
    .A2(_2954_),
    .B1(_2960_),
    .B2(_2961_),
    .C(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7719_ (.A1(_2780_),
    .A2(_2937_),
    .B(_2791_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7720_ (.A1(_2591_),
    .A2(_2963_),
    .B1(_2964_),
    .B2(_2931_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7721_ (.A1(_2775_),
    .A2(_2965_),
    .B(_1471_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7722_ (.A1(_2929_),
    .A2(_2966_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7723_ (.A1(_1644_),
    .A2(_2930_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7724_ (.A1(_1738_),
    .A2(_2967_),
    .Z(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7725_ (.A1(\as2650.pc[6] ),
    .A2(_0723_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7726_ (.I(_2969_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7727_ (.A1(\as2650.pc[5] ),
    .A2(net1),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7728_ (.A1(_2933_),
    .A2(_2971_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7729_ (.A1(_1643_),
    .A2(_0603_),
    .B(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7730_ (.A1(_2886_),
    .A2(_2889_),
    .A3(_2932_),
    .B(_2973_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7731_ (.A1(_2970_),
    .A2(_2974_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7732_ (.A1(_2885_),
    .A2(_2968_),
    .B1(_2975_),
    .B2(_2892_),
    .C(_2758_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7733_ (.A1(_2882_),
    .A2(_2976_),
    .B(_2894_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7734_ (.A1(_2843_),
    .A2(_2975_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7735_ (.A1(_4094_),
    .A2(_2809_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7736_ (.A1(_1374_),
    .A2(_2851_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7737_ (.A1(_2979_),
    .A2(_2980_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7738_ (.A1(_2446_),
    .A2(_2968_),
    .B1(_2981_),
    .B2(_1257_),
    .C(_1317_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7739_ (.A1(_2576_),
    .A2(_2978_),
    .A3(_2982_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7740_ (.A1(_1643_),
    .A2(_1638_),
    .A3(_2907_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7741_ (.A1(_1650_),
    .A2(_2984_),
    .Z(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7742_ (.A1(_0604_),
    .A2(_0531_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7743_ (.I(_0723_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7744_ (.A1(_2987_),
    .A2(_0595_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7745_ (.I(_2988_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7746_ (.A1(_2986_),
    .A2(_2943_),
    .A3(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7747_ (.A1(_2986_),
    .A2(_2943_),
    .B(_2989_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7748_ (.A1(_2546_),
    .A2(_2991_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7749_ (.A1(_1412_),
    .A2(_2868_),
    .B1(_2990_),
    .B2(_2992_),
    .C(_2869_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7750_ (.A1(_2857_),
    .A2(_2985_),
    .B(_2993_),
    .C(_2592_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7751_ (.A1(_2983_),
    .A2(_2994_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7752_ (.I(_2760_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7753_ (.A1(\as2650.stack[4][6] ),
    .A2(_2836_),
    .B1(_1176_),
    .B2(\as2650.stack[5][6] ),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7754_ (.A1(\as2650.stack[7][6] ),
    .A2(_1297_),
    .B1(_2691_),
    .B2(\as2650.stack[6][6] ),
    .C(_0914_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7755_ (.A1(\as2650.stack[3][6] ),
    .A2(_1663_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7756_ (.A1(_0949_),
    .A2(_2999_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7757_ (.A1(\as2650.stack[0][6] ),
    .A2(_2819_),
    .B1(_2694_),
    .B2(\as2650.stack[1][6] ),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7758_ (.I(_3001_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7759_ (.A1(\as2650.stack[2][6] ),
    .A2(_1047_),
    .B(_3000_),
    .C(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7760_ (.A1(_2997_),
    .A2(_2998_),
    .B(_3003_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7761_ (.A1(_2996_),
    .A2(_2968_),
    .B1(_3004_),
    .B2(_2823_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7762_ (.A1(_2976_),
    .A2(_2995_),
    .B(_3005_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7763_ (.A1(_2968_),
    .A2(_2977_),
    .B1(_3006_),
    .B2(_2688_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7764_ (.A1(_1696_),
    .A2(_2878_),
    .B(_2927_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7765_ (.A1(_2830_),
    .A2(_3007_),
    .B(_3008_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7766_ (.A1(_1657_),
    .A2(_2775_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7767_ (.A1(\as2650.pc[6] ),
    .A2(\as2650.pc[5] ),
    .A3(_2930_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7768_ (.A1(_1655_),
    .A2(_3010_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7769_ (.I(\as2650.stack[2][7] ),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7770_ (.A1(\as2650.stack[3][7] ),
    .A2(_1663_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7771_ (.A1(\as2650.stack[0][7] ),
    .A2(_1192_),
    .B1(_2956_),
    .B2(\as2650.stack[1][7] ),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7772_ (.A1(_3012_),
    .A2(_0898_),
    .B1(_3013_),
    .B2(_0912_),
    .C(_3014_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7773_ (.A1(\as2650.stack[7][7] ),
    .A2(_2762_),
    .B1(_1046_),
    .B2(\as2650.stack[6][7] ),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7774_ (.A1(\as2650.stack[4][7] ),
    .A2(_2819_),
    .B1(_2956_),
    .B2(\as2650.stack[5][7] ),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7775_ (.A1(_0922_),
    .A2(_3016_),
    .A3(_3017_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7776_ (.A1(_3015_),
    .A2(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7777_ (.A1(\as2650.pc[7] ),
    .A2(net2),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7778_ (.A1(_1650_),
    .A2(_1373_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7779_ (.A1(_2970_),
    .A2(_2974_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7780_ (.A1(_3021_),
    .A2(_3022_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7781_ (.A1(_3020_),
    .A2(_3023_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7782_ (.A1(_2843_),
    .A2(_3024_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7783_ (.A1(_2599_),
    .A2(_3011_),
    .B(_2489_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7784_ (.A1(_2558_),
    .A2(_2804_),
    .B1(_1430_),
    .B2(_2312_),
    .C(_3026_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7785_ (.A1(_2576_),
    .A2(_3025_),
    .A3(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7786_ (.I(_2704_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7787_ (.A1(_1737_),
    .A2(_2984_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7788_ (.A1(_1794_),
    .A2(_3030_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7789_ (.A1(_1372_),
    .A2(_0595_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7790_ (.A1(net3),
    .A2(_4215_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7791_ (.A1(_3032_),
    .A2(_2991_),
    .B(_3033_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7792_ (.A1(_3032_),
    .A2(_2991_),
    .A3(_3033_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7793_ (.A1(_2897_),
    .A2(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7794_ (.A1(_2558_),
    .A2(_2594_),
    .B1(_3034_),
    .B2(_3036_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7795_ (.A1(_2548_),
    .A2(_2466_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7796_ (.I(_3038_),
    .Z(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7797_ (.I(_2536_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7798_ (.A1(_3029_),
    .A2(_3031_),
    .B1(_3037_),
    .B2(_3039_),
    .C(_3040_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7799_ (.A1(_2892_),
    .A2(_3024_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7800_ (.A1(_2781_),
    .A2(_3011_),
    .B(_2789_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7801_ (.A1(_3028_),
    .A2(_3041_),
    .B(_3042_),
    .C(_3043_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7802_ (.A1(_2832_),
    .A2(_3011_),
    .B1(_3019_),
    .B2(_2842_),
    .C(_3044_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7803_ (.A1(_2779_),
    .A2(_3042_),
    .A3(_3043_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7804_ (.A1(_2438_),
    .A2(_3046_),
    .B(_3011_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7805_ (.A1(_2831_),
    .A2(_3045_),
    .B(_3047_),
    .C(_2829_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7806_ (.I(_2532_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7807_ (.A1(_3009_),
    .A2(_3048_),
    .B(_3049_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7808_ (.I(\as2650.pc[8] ),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7809_ (.I(_3050_),
    .Z(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7810_ (.A1(_1793_),
    .A2(_3010_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7811_ (.A1(_3050_),
    .A2(_3052_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7812_ (.A1(_3050_),
    .A2(_2987_),
    .Z(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7813_ (.A1(_2969_),
    .A2(_3020_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7814_ (.A1(_1794_),
    .A2(_1737_),
    .B(_0724_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7815_ (.A1(_2974_),
    .A2(_3055_),
    .B(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7816_ (.A1(_3054_),
    .A2(_3057_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7817_ (.A1(_2891_),
    .A2(_3058_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7818_ (.A1(_2781_),
    .A2(_3053_),
    .B(_3059_),
    .C(_2789_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7819_ (.A1(_2780_),
    .A2(_3060_),
    .B(_2770_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7820_ (.I(\as2650.addr_buff[0] ),
    .Z(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7821_ (.I(_3062_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7822_ (.A1(_0784_),
    .A2(_4215_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7823_ (.A1(_3064_),
    .A2(_3034_),
    .B(_2320_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7824_ (.A1(_3063_),
    .A2(_3065_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7825_ (.A1(_1088_),
    .A2(_1655_),
    .A3(_3030_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7826_ (.A1(_1656_),
    .A2(_3030_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7827_ (.A1(_3051_),
    .A2(_3068_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7828_ (.A1(_3067_),
    .A2(_3069_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7829_ (.I(_2321_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7830_ (.A1(_3063_),
    .A2(_2861_),
    .B1(_3071_),
    .B2(_1398_),
    .C(_1353_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7831_ (.A1(_1577_),
    .A2(_3053_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7832_ (.A1(_1578_),
    .A2(_3058_),
    .B(_3073_),
    .C(_1248_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7833_ (.A1(_2793_),
    .A2(_3070_),
    .B1(_3072_),
    .B2(_3074_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7834_ (.A1(_2869_),
    .A2(_3066_),
    .B1(_3075_),
    .B2(_2735_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7835_ (.A1(_2592_),
    .A2(_3076_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7836_ (.A1(_2824_),
    .A2(_3053_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7837_ (.A1(_0925_),
    .A2(_2961_),
    .B1(_3060_),
    .B2(_3077_),
    .C(_3078_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7838_ (.A1(_3053_),
    .A2(_3061_),
    .B1(_3079_),
    .B2(_2462_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7839_ (.A1(_2685_),
    .A2(_3080_),
    .B(_2927_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7840_ (.A1(_3051_),
    .A2(_2686_),
    .B(_3081_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7841_ (.I(\as2650.pc[9] ),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7842_ (.I(_3082_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7843_ (.A1(\as2650.pc[9] ),
    .A2(\as2650.pc[8] ),
    .A3(_3052_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7844_ (.A1(_1088_),
    .A2(_3052_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7845_ (.A1(_3083_),
    .A2(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7846_ (.A1(_3084_),
    .A2(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7847_ (.A1(_3082_),
    .A2(_2987_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7848_ (.A1(_1088_),
    .A2(_1371_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7849_ (.A1(_3054_),
    .A2(_3057_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7850_ (.A1(_3089_),
    .A2(_3090_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7851_ (.A1(_3088_),
    .A2(_3091_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7852_ (.A1(_2788_),
    .A2(_3092_),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7853_ (.A1(_2782_),
    .A2(_3087_),
    .B(_3093_),
    .C(_2789_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7854_ (.A1(_3063_),
    .A2(_3065_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7855_ (.A1(_2296_),
    .A2(_3095_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7856_ (.I(\as2650.addr_buff[1] ),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7857_ (.A1(_3097_),
    .A2(_2860_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7858_ (.A1(_2743_),
    .A2(_3098_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7859_ (.A1(_1256_),
    .A2(_3099_),
    .B(_4293_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7860_ (.A1(_2947_),
    .A2(_3092_),
    .B1(_3087_),
    .B2(_2599_),
    .C(_3100_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7861_ (.A1(_1106_),
    .A2(_3067_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7862_ (.A1(_2793_),
    .A2(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7863_ (.A1(_3101_),
    .A2(_3103_),
    .B(_2433_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7864_ (.A1(_3039_),
    .A2(_3096_),
    .B(_3104_),
    .C(_2465_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7865_ (.A1(_0959_),
    .A2(_2961_),
    .B1(_3094_),
    .B2(_3105_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7866_ (.A1(_2779_),
    .A2(_3094_),
    .B(_2996_),
    .C(_2770_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7867_ (.A1(_2732_),
    .A2(_3106_),
    .B1(_3107_),
    .B2(_3087_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7868_ (.A1(_2685_),
    .A2(_3108_),
    .B(_2927_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7869_ (.A1(_3083_),
    .A2(_2686_),
    .B(_3109_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7870_ (.A1(_1114_),
    .A2(_2775_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7871_ (.I(\as2650.pc[10] ),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7872_ (.A1(_3111_),
    .A2(_3084_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7873_ (.I(_3112_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7874_ (.A1(_3062_),
    .A2(_3097_),
    .A3(_3065_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7875_ (.A1(_2298_),
    .A2(_3114_),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7876_ (.A1(_3083_),
    .A2(_3067_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7877_ (.A1(_3111_),
    .A2(_3116_),
    .Z(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7878_ (.A1(\as2650.pc[10] ),
    .A2(_2987_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7879_ (.I(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7880_ (.I(_3119_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7881_ (.A1(_3090_),
    .A2(_3088_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7882_ (.A1(\as2650.pc[9] ),
    .A2(_1371_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7883_ (.A1(_3089_),
    .A2(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7884_ (.A1(_3121_),
    .A2(_3123_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7885_ (.A1(_3120_),
    .A2(_3124_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7886_ (.A1(\as2650.addr_buff[2] ),
    .A2(_0290_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7887_ (.A1(_0349_),
    .A2(_2260_),
    .B(_3126_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7888_ (.A1(_1255_),
    .A2(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7889_ (.A1(_1797_),
    .A2(_3128_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7890_ (.A1(_2843_),
    .A2(_3125_),
    .B1(_3112_),
    .B2(_2796_),
    .C(_3129_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _7891_ (.A1(_3039_),
    .A2(_3115_),
    .B1(_3117_),
    .B2(_3029_),
    .C1(_2600_),
    .C2(_3130_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7892_ (.A1(_2891_),
    .A2(_3125_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7893_ (.A1(_2781_),
    .A2(_3113_),
    .B(_3132_),
    .C(_2335_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7894_ (.A1(_2470_),
    .A2(_3131_),
    .B(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7895_ (.A1(_0980_),
    .A2(_2842_),
    .B1(_3113_),
    .B2(_2832_),
    .C(_3134_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7896_ (.A1(_2779_),
    .A2(_3133_),
    .B(_2770_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7897_ (.A1(_3113_),
    .A2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7898_ (.A1(_2831_),
    .A2(_3135_),
    .B(_3137_),
    .C(_2829_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7899_ (.A1(_3110_),
    .A2(_3138_),
    .B(_3049_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7900_ (.I(\as2650.pc[11] ),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7901_ (.A1(_3111_),
    .A2(_3084_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7902_ (.I(_3140_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7903_ (.A1(_3139_),
    .A2(_3141_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7904_ (.I(\as2650.addr_buff[3] ),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7905_ (.A1(\as2650.addr_buff[0] ),
    .A2(_3097_),
    .A3(\as2650.addr_buff[2] ),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7906_ (.A1(_3064_),
    .A2(_3034_),
    .B(_3144_),
    .C(_2545_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7907_ (.A1(_3143_),
    .A2(_3145_),
    .Z(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7908_ (.A1(\as2650.pc[11] ),
    .A2(_0726_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7909_ (.A1(\as2650.pc[10] ),
    .A2(_1491_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7910_ (.A1(_3120_),
    .A2(_3124_),
    .B(_3148_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7911_ (.A1(_3147_),
    .A2(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7912_ (.A1(_3143_),
    .A2(_2803_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7913_ (.A1(_0431_),
    .A2(_2593_),
    .B(_2354_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7914_ (.A1(_2796_),
    .A2(_3142_),
    .B1(_3151_),
    .B2(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7915_ (.A1(_2947_),
    .A2(_3150_),
    .B(_3153_),
    .C(_1285_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7916_ (.A1(_3111_),
    .A2(_3083_),
    .A3(_3067_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7917_ (.A1(_1121_),
    .A2(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7918_ (.A1(_3139_),
    .A2(_3141_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7919_ (.A1(_2736_),
    .A2(_3157_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7920_ (.A1(_2736_),
    .A2(_3156_),
    .B(_3158_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7921_ (.A1(_2280_),
    .A2(_3159_),
    .B(_2735_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7922_ (.A1(_2472_),
    .A2(_3150_),
    .B1(_3157_),
    .B2(_2647_),
    .C(_2537_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7923_ (.A1(_2706_),
    .A2(_3142_),
    .B1(_3154_),
    .B2(_3160_),
    .C(_3161_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7924_ (.A1(_2813_),
    .A2(_3146_),
    .B(_3162_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7925_ (.A1(_0994_),
    .A2(_2690_),
    .B1(_3157_),
    .B2(_2689_),
    .C(_2687_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7926_ (.A1(_2894_),
    .A2(_3142_),
    .B1(_3163_),
    .B2(_3164_),
    .C(_2684_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7927_ (.A1(_1122_),
    .A2(_2686_),
    .B(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7928_ (.A1(_2640_),
    .A2(_3166_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7929_ (.A1(_1120_),
    .A2(_3141_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7930_ (.A1(_1129_),
    .A2(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7931_ (.A1(_3119_),
    .A2(_3147_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7932_ (.A1(_1120_),
    .A2(_1491_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7933_ (.A1(_3089_),
    .A2(_3122_),
    .A3(_3148_),
    .A4(_3170_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7934_ (.A1(_3121_),
    .A2(_3169_),
    .B(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7935_ (.A1(_1128_),
    .A2(_1373_),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7936_ (.A1(_3172_),
    .A2(_3173_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7937_ (.A1(_2788_),
    .A2(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7938_ (.A1(_2885_),
    .A2(_3168_),
    .B(_3175_),
    .C(_2758_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7939_ (.A1(_2882_),
    .A2(_3176_),
    .B(_2894_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7940_ (.A1(_3143_),
    .A2(_3145_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7941_ (.A1(_2306_),
    .A2(_3178_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7942_ (.A1(\as2650.addr_buff[4] ),
    .A2(_2803_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7943_ (.A1(_2905_),
    .A2(_3180_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7944_ (.A1(_2796_),
    .A2(_3168_),
    .B1(_3181_),
    .B2(_1256_),
    .C(_1354_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7945_ (.A1(_2947_),
    .A2(_3174_),
    .B(_3182_),
    .C(_2600_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7946_ (.A1(_1121_),
    .A2(_3155_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7947_ (.A1(_1129_),
    .A2(_3184_),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7948_ (.A1(_3029_),
    .A2(_3185_),
    .B(_2465_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7949_ (.A1(_2813_),
    .A2(_3179_),
    .B(_3183_),
    .C(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7950_ (.A1(_2760_),
    .A2(_3168_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7951_ (.A1(_1008_),
    .A2(_2842_),
    .B1(_3176_),
    .B2(_3187_),
    .C(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7952_ (.A1(_3168_),
    .A2(_3177_),
    .B1(_3189_),
    .B2(_2688_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7953_ (.I(_2338_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7954_ (.A1(_1130_),
    .A2(_2829_),
    .B(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7955_ (.A1(_2830_),
    .A2(_3190_),
    .B(_3192_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7956_ (.A1(_1128_),
    .A2(_3139_),
    .A3(_3141_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7957_ (.A1(_1135_),
    .A2(_3193_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7958_ (.A1(_2306_),
    .A2(_3178_),
    .B(_2948_),
    .C(_3039_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7959_ (.A1(_1129_),
    .A2(_1121_),
    .A3(_3155_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7960_ (.A1(_1135_),
    .A2(_3196_),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7961_ (.A1(_4095_),
    .A2(_2861_),
    .B(_2708_),
    .C(_1353_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7962_ (.A1(_2599_),
    .A2(_3194_),
    .B(_3198_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7963_ (.A1(_2537_),
    .A2(_3199_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7964_ (.A1(_2857_),
    .A2(_3197_),
    .B1(_3194_),
    .B2(_2882_),
    .C(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7965_ (.A1(_3195_),
    .A2(_3201_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7966_ (.A1(_1021_),
    .A2(_2961_),
    .B1(_3194_),
    .B2(_2996_),
    .C(_3202_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7967_ (.A1(_2462_),
    .A2(_2782_),
    .B(_3194_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7968_ (.A1(_2591_),
    .A2(_3203_),
    .B(_3204_),
    .C(_2685_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7969_ (.A1(_1135_),
    .A2(_2731_),
    .B(_2339_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7970_ (.A1(_3205_),
    .A2(_3206_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7971_ (.A1(\as2650.pc[13] ),
    .A2(\as2650.pc[12] ),
    .A3(_1120_),
    .A4(_3140_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7972_ (.A1(\as2650.pc[14] ),
    .A2(_3207_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7973_ (.A1(_2462_),
    .A2(_3208_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7974_ (.A1(\as2650.pc[13] ),
    .A2(_1128_),
    .A3(_3139_),
    .A4(_3155_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7975_ (.A1(\as2650.pc[14] ),
    .A2(_3210_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7976_ (.A1(_3038_),
    .A2(_2979_),
    .B1(_3211_),
    .B2(_3029_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7977_ (.A1(_4094_),
    .A2(_2861_),
    .B1(_2445_),
    .B2(_3208_),
    .C(_2433_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7978_ (.A1(_2464_),
    .A2(_3213_),
    .B(_1335_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7979_ (.A1(_1548_),
    .A2(_3212_),
    .B(_3214_),
    .C(_2335_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7980_ (.A1(_2701_),
    .A2(_2778_),
    .B(_3208_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7981_ (.A1(_2461_),
    .A2(_3215_),
    .B(_3216_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7982_ (.A1(_1034_),
    .A2(_2690_),
    .B1(_3208_),
    .B2(_2689_),
    .C(_3217_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7983_ (.A1(_3209_),
    .A2(_3218_),
    .B(_2727_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7984_ (.A1(\as2650.pc[14] ),
    .A2(_2731_),
    .B(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7985_ (.A1(_2640_),
    .A2(_3220_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7986_ (.A1(_2268_),
    .A2(_4081_),
    .A3(_2393_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7987_ (.A1(_2530_),
    .A2(_2406_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7988_ (.A1(_2331_),
    .A2(_3221_),
    .A3(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7989_ (.A1(_1243_),
    .A2(_1352_),
    .A3(_2656_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7990_ (.A1(_1567_),
    .A2(_2417_),
    .A3(_3224_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7991_ (.A1(_2561_),
    .A2(_4262_),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7992_ (.A1(_4363_),
    .A2(_3226_),
    .B(_4260_),
    .C(_2656_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7993_ (.A1(_2652_),
    .A2(_2673_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7994_ (.A1(_4133_),
    .A2(_2676_),
    .A3(_2276_),
    .A4(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7995_ (.A1(_1093_),
    .A2(_1437_),
    .A3(_3227_),
    .A4(_3229_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7996_ (.A1(_1434_),
    .A2(_2400_),
    .A3(_3225_),
    .A4(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7997_ (.A1(_2860_),
    .A2(_4396_),
    .B1(_1843_),
    .B2(_4096_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7998_ (.A1(_4364_),
    .A2(_4060_),
    .A3(_1431_),
    .B1(_3232_),
    .B2(_2268_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7999_ (.A1(_1443_),
    .A2(_2562_),
    .B(_1343_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8000_ (.A1(_1078_),
    .A2(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8001_ (.A1(_1420_),
    .A2(_3235_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8002_ (.A1(_1467_),
    .A2(_3231_),
    .A3(_3233_),
    .A4(_3236_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8003_ (.A1(_1271_),
    .A2(_1352_),
    .A3(_0352_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8004_ (.A1(_4079_),
    .A2(_1433_),
    .B(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8005_ (.A1(_1345_),
    .A2(_1455_),
    .B1(_3239_),
    .B2(_2656_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8006_ (.A1(_2422_),
    .A2(_3240_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8007_ (.A1(_3223_),
    .A2(_3237_),
    .A3(_3241_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8008_ (.I(_3242_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8009_ (.I(_3243_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8010_ (.I(_3244_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8011_ (.I(_2377_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8012_ (.A1(_4004_),
    .A2(_1218_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8013_ (.I(_3247_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8014_ (.I(_3248_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8015_ (.A1(\as2650.carry ),
    .A2(_3249_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8016_ (.A1(_4005_),
    .A2(_1219_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8017_ (.I(_3251_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8018_ (.I(_0887_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8019_ (.A1(_0905_),
    .A2(_3252_),
    .B(_3253_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8020_ (.A1(_0880_),
    .A2(_2700_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8021_ (.A1(_3250_),
    .A2(_3254_),
    .B(_3246_),
    .C(_3255_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8022_ (.A1(_4322_),
    .A2(_3246_),
    .B(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8023_ (.I(_1387_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8024_ (.I(_2349_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8025_ (.A1(_1383_),
    .A2(_3258_),
    .B1(_4224_),
    .B2(_1528_),
    .C(_3259_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8026_ (.A1(_1422_),
    .A2(_3257_),
    .B(_3260_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8027_ (.I(_4379_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8028_ (.I(_1462_),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8029_ (.I(_1464_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8030_ (.A1(_3262_),
    .A2(_3263_),
    .B1(_3264_),
    .B2(_1559_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8031_ (.A1(_1580_),
    .A2(_4250_),
    .B(_3265_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8032_ (.A1(_3244_),
    .A2(_3261_),
    .A3(_3266_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8033_ (.I(_2547_),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8034_ (.I(_1426_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8035_ (.I(_3269_),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8036_ (.I(_2626_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8037_ (.A1(_3271_),
    .A2(_4272_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8038_ (.I(_2898_),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8039_ (.A1(_3271_),
    .A2(_4279_),
    .B(_3272_),
    .C(_3273_),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8040_ (.A1(_3268_),
    .A2(_4186_),
    .B(_3270_),
    .C(_3274_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8041_ (.A1(_1709_),
    .A2(_3245_),
    .B1(_3267_),
    .B2(_3275_),
    .C(_2590_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8042_ (.I(_3243_),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8043_ (.I(_2622_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8044_ (.A1(_3277_),
    .A2(_4359_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8045_ (.A1(_3277_),
    .A2(_4374_),
    .B(_3278_),
    .C(_3273_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8046_ (.A1(_3268_),
    .A2(_4355_),
    .B(_3270_),
    .C(_3279_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8047_ (.I(_1267_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8048_ (.I(_0934_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8049_ (.I(_3247_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8050_ (.A1(_0902_),
    .A2(_3283_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8051_ (.A1(_1511_),
    .A2(_3283_),
    .B(_3284_),
    .C(_0886_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8052_ (.A1(_0887_),
    .A2(_2767_),
    .B(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8053_ (.A1(_4417_),
    .A2(_0934_),
    .B(_4078_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8054_ (.A1(_3282_),
    .A2(_3286_),
    .B(_3287_),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8055_ (.A1(_1381_),
    .A2(_3262_),
    .B(_3288_),
    .C(_1267_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8056_ (.A1(_3281_),
    .A2(_0355_),
    .B(_3289_),
    .C(_1395_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8057_ (.A1(_1401_),
    .A2(_1396_),
    .B(_3290_),
    .C(_2603_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8058_ (.A1(_2336_),
    .A2(_4400_),
    .B(_3291_),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8059_ (.A1(_3258_),
    .A2(_2651_),
    .B1(_3292_),
    .B2(_1474_),
    .C(_3243_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8060_ (.A1(_1721_),
    .A2(_3276_),
    .B1(_3280_),
    .B2(_3293_),
    .C(_2639_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8061_ (.I(_3269_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8062_ (.A1(_2256_),
    .A2(_0327_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8063_ (.A1(_2623_),
    .A2(_0331_),
    .B(_3295_),
    .C(_2547_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8064_ (.A1(_3273_),
    .A2(_0316_),
    .B(_3294_),
    .C(_3296_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8065_ (.A1(\as2650.overflow ),
    .A2(_3249_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8066_ (.A1(_1173_),
    .A2(_3252_),
    .B(_0936_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8067_ (.A1(_0879_),
    .A2(_2822_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8068_ (.A1(_3298_),
    .A2(_3299_),
    .B(_0935_),
    .C(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8069_ (.A1(_0370_),
    .A2(_3246_),
    .B(_3301_),
    .C(_1527_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8070_ (.I(_1365_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8071_ (.A1(_3303_),
    .A2(_3258_),
    .B(_1385_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8072_ (.A1(_1385_),
    .A2(_1495_),
    .B1(_3302_),
    .B2(_3304_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8073_ (.A1(_2299_),
    .A2(_3264_),
    .B1(_3259_),
    .B2(_3305_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8074_ (.A1(_1568_),
    .A2(_0357_),
    .B1(_3263_),
    .B2(_2014_),
    .C(_3243_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8075_ (.A1(_3297_),
    .A2(_3306_),
    .A3(_3307_),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8076_ (.A1(_1619_),
    .A2(_3245_),
    .B(_3308_),
    .C(_2730_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8077_ (.A1(_3271_),
    .A2(_0452_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8078_ (.A1(_3277_),
    .A2(_0458_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8079_ (.A1(_3268_),
    .A2(_3309_),
    .A3(_3310_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8080_ (.A1(_3268_),
    .A2(_0413_),
    .B(_3270_),
    .C(_3311_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8081_ (.I(_3281_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8082_ (.A1(_4206_),
    .A2(_3249_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8083_ (.A1(\as2650.psu[3] ),
    .A2(_3252_),
    .B(_0936_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8084_ (.A1(_3253_),
    .A2(_2841_),
    .B1(_3314_),
    .B2(_3315_),
    .C(_0935_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8085_ (.A1(_0470_),
    .A2(_3246_),
    .B(_3316_),
    .C(_1528_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8086_ (.A1(_3303_),
    .A2(_2014_),
    .B(_1385_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8087_ (.A1(_3313_),
    .A2(_0428_),
    .B1(_3317_),
    .B2(_3318_),
    .ZN(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8088_ (.A1(_1388_),
    .A2(_2494_),
    .B(_3242_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8089_ (.A1(_1580_),
    .A2(_0436_),
    .B(_3320_),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8090_ (.A1(_2303_),
    .A2(_3264_),
    .B1(_3259_),
    .B2(_3319_),
    .C(_3321_),
    .ZN(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8091_ (.A1(_1628_),
    .A2(_3276_),
    .B1(_3312_),
    .B2(_3322_),
    .C(_2639_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8092_ (.A1(_3277_),
    .A2(_0553_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8093_ (.I(_2594_),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8094_ (.A1(_3271_),
    .A2(_0516_),
    .B(_3324_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8095_ (.I(_2261_),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8096_ (.A1(_3326_),
    .A2(_0510_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8097_ (.A1(_3323_),
    .A2(_3325_),
    .B(_3270_),
    .C(_3327_),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8098_ (.A1(_4286_),
    .A2(_3251_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8099_ (.A1(_1490_),
    .A2(_3252_),
    .B(_3329_),
    .C(_0936_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8100_ (.A1(_3253_),
    .A2(_2923_),
    .B(_3330_),
    .C(_0935_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8101_ (.A1(_1951_),
    .A2(_0873_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8102_ (.A1(_1422_),
    .A2(_3331_),
    .A3(_3332_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8103_ (.A1(_1381_),
    .A2(_1495_),
    .B1(_0714_),
    .B2(_3281_),
    .C(_1395_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8104_ (.A1(_1411_),
    .A2(_1395_),
    .B1(_3333_),
    .B2(_3334_),
    .C(_2586_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8105_ (.A1(_1569_),
    .A2(_0543_),
    .B1(_2651_),
    .B2(_0428_),
    .C(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8106_ (.A1(_3328_),
    .A2(_3336_),
    .B(_3276_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8107_ (.A1(_2177_),
    .A2(_3245_),
    .B(_3337_),
    .C(_2730_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8108_ (.I(_2532_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8109_ (.A1(_3324_),
    .A2(_2096_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8110_ (.I(_2626_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8111_ (.A1(_3340_),
    .A2(_0619_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8112_ (.A1(_2623_),
    .A2(_0587_),
    .B(_2547_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8113_ (.A1(_3341_),
    .A2(_3342_),
    .B(_3269_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8114_ (.A1(_1365_),
    .A2(_0591_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8115_ (.A1(\as2650.psu[5] ),
    .A2(_3251_),
    .ZN(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8116_ (.A1(\as2650.psl[5] ),
    .A2(_3248_),
    .B(_0886_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8117_ (.A1(_0875_),
    .A2(_2960_),
    .ZN(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8118_ (.A1(_3345_),
    .A2(_3346_),
    .B(_3347_),
    .C(_3282_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8119_ (.A1(_0526_),
    .A2(_2377_),
    .B(_3348_),
    .C(_1527_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8120_ (.A1(_3344_),
    .A2(_3349_),
    .B(_3281_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8121_ (.A1(_1479_),
    .A2(_1386_),
    .B(_4101_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8122_ (.A1(_1287_),
    .A2(_1363_),
    .B1(_3350_),
    .B2(_3351_),
    .C(_2724_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8123_ (.A1(_2431_),
    .A2(_0607_),
    .B(_3352_),
    .C(_1473_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8124_ (.A1(_0714_),
    .A2(_3263_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8125_ (.A1(_3339_),
    .A2(_3343_),
    .B(_3353_),
    .C(_3354_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8126_ (.I0(_3355_),
    .I1(_1734_),
    .S(_3244_),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8127_ (.A1(_3338_),
    .A2(_3356_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8128_ (.A1(_2482_),
    .A2(_0709_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8129_ (.A1(_3340_),
    .A2(_0735_),
    .B(_2898_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8130_ (.A1(_3324_),
    .A2(_0700_),
    .B1(_3357_),
    .B2(_3358_),
    .C(_3269_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8131_ (.A1(_1375_),
    .A2(_3248_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8132_ (.A1(_1492_),
    .A2(_3248_),
    .B(_3360_),
    .C(_0879_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8133_ (.A1(_0880_),
    .A2(_3004_),
    .B(_3361_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8134_ (.A1(_2036_),
    .A2(_0873_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8135_ (.A1(_0873_),
    .A2(_3362_),
    .B(_3363_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8136_ (.A1(_1479_),
    .A2(_4223_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8137_ (.A1(_1381_),
    .A2(_0646_),
    .B1(_3364_),
    .B2(_1422_),
    .C(_3365_),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8138_ (.A1(_1386_),
    .A2(_3263_),
    .B1(_3259_),
    .B2(_3366_),
    .C1(_3264_),
    .C2(_0726_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8139_ (.A1(_1580_),
    .A2(_0721_),
    .B(_3359_),
    .C(_3367_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8140_ (.I0(_3368_),
    .I1(_0713_),
    .S(_3244_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8141_ (.A1(_3338_),
    .A2(_3369_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8142_ (.A1(_2623_),
    .A2(_0781_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8143_ (.A1(_3340_),
    .A2(_0797_),
    .B(_3324_),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _8144_ (.A1(_3273_),
    .A2(_1475_),
    .B1(_3370_),
    .B2(_3371_),
    .C(_3294_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8145_ (.A1(_1487_),
    .A2(_3283_),
    .B(_0875_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8146_ (.A1(_1518_),
    .A2(_3283_),
    .B(_3373_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8147_ (.A1(_0887_),
    .A2(_3019_),
    .B(_3374_),
    .C(_3282_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8148_ (.A1(_2076_),
    .A2(_2377_),
    .B(_3375_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8149_ (.A1(_1527_),
    .A2(_3376_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8150_ (.A1(_1479_),
    .A2(_1366_),
    .A3(_3377_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8151_ (.A1(_1480_),
    .A2(_3378_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8152_ (.A1(_1363_),
    .A2(_3379_),
    .B(_2586_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8153_ (.A1(_1569_),
    .A2(_0787_),
    .B1(_1397_),
    .B2(_3380_),
    .C1(_2651_),
    .C2(_1340_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8154_ (.A1(_3372_),
    .A2(_3381_),
    .B(_3276_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8155_ (.A1(_1653_),
    .A2(_3245_),
    .B(_3382_),
    .C(_2730_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8156_ (.A1(_1173_),
    .A2(_0920_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8157_ (.A1(_1592_),
    .A2(_3383_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8158_ (.I(_3384_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8159_ (.I(_3385_),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8160_ (.A1(_1602_),
    .A2(_1160_),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8161_ (.I(_3387_),
    .Z(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8162_ (.A1(_1747_),
    .A2(_0973_),
    .A3(_1750_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8163_ (.I(_3389_),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8164_ (.A1(_1598_),
    .A2(_3388_),
    .B1(_3390_),
    .B2(\as2650.stack[6][0] ),
    .C(_3385_),
    .ZN(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8165_ (.A1(_1709_),
    .A2(_3386_),
    .B(_3391_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8166_ (.A1(_1614_),
    .A2(_3388_),
    .B1(_3390_),
    .B2(\as2650.stack[6][1] ),
    .C(_3384_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8167_ (.A1(_1721_),
    .A2(_3386_),
    .B(_3392_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8168_ (.I(_3389_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8169_ (.A1(\as2650.stack[6][2] ),
    .A2(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8170_ (.I(_3387_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8171_ (.I(_3384_),
    .Z(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8172_ (.A1(_1679_),
    .A2(_3395_),
    .B(_3396_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8173_ (.A1(_1675_),
    .A2(_3386_),
    .B1(_3394_),
    .B2(_3397_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8174_ (.I(_3385_),
    .Z(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8175_ (.A1(\as2650.stack[6][3] ),
    .A2(_3393_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8176_ (.A1(_1729_),
    .A2(_3395_),
    .B(_3396_),
    .ZN(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8177_ (.A1(_1727_),
    .A2(_3398_),
    .B1(_3399_),
    .B2(_3400_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8178_ (.A1(\as2650.stack[6][4] ),
    .A2(_3393_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8179_ (.A1(_1640_),
    .A2(_3395_),
    .B(_3396_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8180_ (.A1(_2177_),
    .A2(_3398_),
    .B1(_3401_),
    .B2(_3402_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8181_ (.A1(\as2650.stack[6][5] ),
    .A2(_3393_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8182_ (.A1(_1693_),
    .A2(_3395_),
    .B(_3396_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8183_ (.A1(_1734_),
    .A2(_3398_),
    .B1(_3403_),
    .B2(_3404_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8184_ (.A1(\as2650.stack[6][6] ),
    .A2(_3390_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8185_ (.A1(_1696_),
    .A2(_3388_),
    .B(_3385_),
    .ZN(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8186_ (.A1(_1648_),
    .A2(_3398_),
    .B1(_3405_),
    .B2(_3406_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8187_ (.A1(_1741_),
    .A2(_3388_),
    .B1(_3390_),
    .B2(\as2650.stack[6][7] ),
    .C(_3384_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8188_ (.A1(_1698_),
    .A2(_3386_),
    .B(_3407_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8189_ (.A1(_1174_),
    .A2(_1298_),
    .A3(_1591_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8190_ (.I(_3408_),
    .Z(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8191_ (.I(_3409_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8192_ (.A1(_1146_),
    .A2(_0900_),
    .A3(_1605_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8193_ (.I(_3411_),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8194_ (.I(_3412_),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8195_ (.A1(\as2650.stack[7][0] ),
    .A2(_3413_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8196_ (.A1(_1602_),
    .A2(_3383_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8197_ (.I(_3415_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8198_ (.I(_3408_),
    .Z(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8199_ (.A1(_1599_),
    .A2(_3416_),
    .B(_3417_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8200_ (.A1(_1709_),
    .A2(_3410_),
    .B1(_3414_),
    .B2(_3418_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8201_ (.I(_3409_),
    .Z(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8202_ (.A1(\as2650.stack[7][1] ),
    .A2(_3412_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8203_ (.A1(_1670_),
    .A2(_3415_),
    .B(_3420_),
    .C(_3409_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8204_ (.A1(_1721_),
    .A2(_3419_),
    .B(_3421_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8205_ (.A1(\as2650.stack[7][2] ),
    .A2(_3413_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8206_ (.A1(_1624_),
    .A2(_3416_),
    .B(_3417_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8207_ (.A1(_1675_),
    .A2(_3410_),
    .B1(_3422_),
    .B2(_3423_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8208_ (.I(_3411_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8209_ (.A1(_1684_),
    .A2(_3424_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8210_ (.A1(\as2650.stack[7][3] ),
    .A2(_3424_),
    .B(_3425_),
    .C(_3409_),
    .ZN(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8211_ (.A1(_1727_),
    .A2(_3419_),
    .B(_3426_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8212_ (.A1(\as2650.stack[7][4] ),
    .A2(_3413_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8213_ (.A1(_1640_),
    .A2(_3416_),
    .B(_3417_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8214_ (.A1(_2177_),
    .A2(_3410_),
    .B1(_3427_),
    .B2(_3428_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8215_ (.A1(\as2650.stack[7][5] ),
    .A2(_3413_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8216_ (.A1(_1646_),
    .A2(_3416_),
    .B(_3417_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8217_ (.A1(_1734_),
    .A2(_3410_),
    .B1(_3429_),
    .B2(_3430_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8218_ (.A1(_1738_),
    .A2(_3412_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8219_ (.A1(\as2650.stack[7][6] ),
    .A2(_3424_),
    .B(_3431_),
    .C(_3408_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8220_ (.A1(_1648_),
    .A2(_3419_),
    .B(_3432_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8221_ (.A1(_1794_),
    .A2(_3412_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8222_ (.A1(\as2650.stack[7][7] ),
    .A2(_3424_),
    .B(_3433_),
    .C(_3408_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8223_ (.A1(_1698_),
    .A2(_3419_),
    .B(_3434_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8224_ (.A1(_1145_),
    .A2(_3383_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8225_ (.I(_3435_),
    .Z(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8226_ (.I(_3436_),
    .Z(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8227_ (.I(_3436_),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8228_ (.A1(\as2650.stack[7][8] ),
    .A2(_3438_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8229_ (.A1(_1190_),
    .A2(_3437_),
    .B(_3439_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8230_ (.I(_3435_),
    .Z(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8231_ (.A1(\as2650.stack[7][9] ),
    .A2(_3440_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8232_ (.A1(_1200_),
    .A2(_3437_),
    .B(_3441_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8233_ (.A1(\as2650.stack[7][10] ),
    .A2(_3440_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8234_ (.A1(_1203_),
    .A2(_3437_),
    .B(_3442_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8235_ (.A1(\as2650.stack[7][11] ),
    .A2(_3440_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8236_ (.A1(_1205_),
    .A2(_3437_),
    .B(_3443_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8237_ (.A1(\as2650.stack[7][12] ),
    .A2(_3440_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8238_ (.A1(_1207_),
    .A2(_3438_),
    .B(_3444_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8239_ (.A1(\as2650.stack[7][13] ),
    .A2(_3436_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8240_ (.A1(_1209_),
    .A2(_3438_),
    .B(_3445_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8241_ (.A1(\as2650.stack[7][14] ),
    .A2(_3436_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8242_ (.A1(_1211_),
    .A2(_3438_),
    .B(_3446_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8243_ (.I(net28),
    .Z(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8244_ (.A1(_2675_),
    .A2(_1561_),
    .B(_2665_),
    .C(_1050_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8245_ (.A1(_2402_),
    .A2(_3448_),
    .ZN(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8246_ (.A1(_2419_),
    .A2(_2423_),
    .A3(_3449_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8247_ (.A1(_1064_),
    .A2(_2394_),
    .B(_2330_),
    .C(_1437_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8248_ (.A1(_2258_),
    .A2(_2382_),
    .B(_3451_),
    .C(_2264_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8249_ (.A1(_2375_),
    .A2(_2666_),
    .A3(_3450_),
    .A4(_3452_),
    .ZN(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8250_ (.A1(_2284_),
    .A2(_2266_),
    .B(_1562_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8251_ (.A1(_2311_),
    .A2(_1442_),
    .A3(_2416_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8252_ (.A1(_3454_),
    .A2(_3455_),
    .B(_1334_),
    .C(_2883_),
    .ZN(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8253_ (.A1(_2399_),
    .A2(_3453_),
    .A3(_3456_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8254_ (.A1(_2391_),
    .A2(_3457_),
    .ZN(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8255_ (.I(_3458_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8256_ (.I(_3459_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8257_ (.I(_2571_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8258_ (.A1(_2620_),
    .A2(_2713_),
    .ZN(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8259_ (.I(_2405_),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8260_ (.I(_2287_),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8261_ (.I(_4365_),
    .Z(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8262_ (.A1(_3465_),
    .A2(_4279_),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8263_ (.A1(_1398_),
    .A2(_3466_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8264_ (.I(_4262_),
    .Z(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8265_ (.A1(_3468_),
    .A2(_4272_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8266_ (.A1(_1496_),
    .A2(_3469_),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8267_ (.A1(_3464_),
    .A2(_3467_),
    .B1(_3470_),
    .B2(_2256_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8268_ (.I(_2272_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8269_ (.A1(_2267_),
    .A2(_2489_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8270_ (.A1(_3447_),
    .A2(_3463_),
    .B1(_3471_),
    .B2(_3472_),
    .C(_3473_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8271_ (.A1(_2606_),
    .A2(_2469_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8272_ (.A1(_1398_),
    .A2(_2897_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8273_ (.A1(_3447_),
    .A2(_2546_),
    .B(_3476_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8274_ (.A1(_2701_),
    .A2(_2713_),
    .B1(_3475_),
    .B2(_3477_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8275_ (.A1(_1553_),
    .A2(_1547_),
    .B(_2471_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8276_ (.I(_3479_),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8277_ (.A1(_2473_),
    .A2(_3478_),
    .B1(_3480_),
    .B2(_1667_),
    .ZN(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8278_ (.A1(_3462_),
    .A2(_3474_),
    .B1(_3481_),
    .B2(_1473_),
    .ZN(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8279_ (.A1(_2494_),
    .A2(_2571_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8280_ (.I(_3483_),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8281_ (.I(_3458_),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8282_ (.A1(_3461_),
    .A2(_3482_),
    .B1(_3484_),
    .B2(_1765_),
    .C(_3485_),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8283_ (.A1(_3447_),
    .A2(_3460_),
    .B(_3486_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8284_ (.A1(_3338_),
    .A2(_3487_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8285_ (.I(_3459_),
    .Z(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8286_ (.I(_3488_),
    .Z(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8287_ (.I(_3483_),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8288_ (.I(_3479_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8289_ (.A1(_1248_),
    .A2(_1547_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8290_ (.I(_3492_),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8291_ (.A1(net53),
    .A2(_3447_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8292_ (.A1(_2804_),
    .A2(_3494_),
    .B(_2750_),
    .ZN(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8293_ (.A1(_3040_),
    .A2(_2749_),
    .B1(_3493_),
    .B2(_3495_),
    .ZN(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8294_ (.I(_3496_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8295_ (.I(_2472_),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8296_ (.A1(_1613_),
    .A2(_3491_),
    .B1(_3497_),
    .B2(_3498_),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8297_ (.I(_2559_),
    .Z(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8298_ (.A1(_2712_),
    .A2(_2748_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8299_ (.A1(_1496_),
    .A2(_4278_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8300_ (.A1(_4393_),
    .A2(_4359_),
    .A3(_3502_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8301_ (.A1(_1400_),
    .A2(_3465_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8302_ (.A1(_2269_),
    .A2(_2270_),
    .A3(_2271_),
    .ZN(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8303_ (.A1(_4090_),
    .A2(_3505_),
    .ZN(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8304_ (.A1(_2625_),
    .A2(_3506_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8305_ (.A1(_3465_),
    .A2(_3503_),
    .B(_3504_),
    .C(_3507_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8306_ (.I(_3468_),
    .Z(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8307_ (.A1(_4241_),
    .A2(_4271_),
    .ZN(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8308_ (.A1(_4391_),
    .A2(_4373_),
    .Z(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8309_ (.A1(_3510_),
    .A2(_3511_),
    .Z(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8310_ (.A1(_3468_),
    .A2(_3512_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8311_ (.A1(_1502_),
    .A2(_3509_),
    .B(_3513_),
    .C(_2625_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8312_ (.I(_2403_),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8313_ (.A1(_3508_),
    .A2(_3514_),
    .B(_3515_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8314_ (.I(_2409_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8315_ (.A1(_3463_),
    .A2(_3494_),
    .B(_3516_),
    .C(_3517_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8316_ (.I(_3473_),
    .Z(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8317_ (.A1(_3500_),
    .A2(_3501_),
    .B(_3518_),
    .C(_3519_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8318_ (.A1(_1360_),
    .A2(_3499_),
    .B(_3520_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8319_ (.A1(_1615_),
    .A2(_3490_),
    .B1(_3521_),
    .B2(_2572_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8320_ (.I(_3459_),
    .Z(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8321_ (.A1(net29),
    .A2(_3523_),
    .B(_3191_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8322_ (.A1(_3489_),
    .A2(_3522_),
    .B(_3524_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8323_ (.I(_3479_),
    .Z(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8324_ (.A1(net53),
    .A2(net28),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8325_ (.A1(net30),
    .A2(_3526_),
    .Z(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8326_ (.A1(_2803_),
    .A2(_3527_),
    .ZN(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8327_ (.A1(_1405_),
    .A2(_2261_),
    .B(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8328_ (.A1(_2884_),
    .A2(_2787_),
    .B1(_3475_),
    .B2(_3529_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8329_ (.A1(_1622_),
    .A2(_3525_),
    .B1(_3530_),
    .B2(_2473_),
    .ZN(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8330_ (.I(_3531_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8331_ (.A1(\as2650.pc[0] ),
    .A2(net5),
    .B(_2748_),
    .ZN(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8332_ (.A1(_2783_),
    .A2(_3533_),
    .B(_2786_),
    .ZN(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8333_ (.A1(_2783_),
    .A2(_2786_),
    .A3(_3533_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8334_ (.A1(_3517_),
    .A2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8335_ (.I(_3505_),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8336_ (.A1(_4391_),
    .A2(_4358_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8337_ (.A1(_4392_),
    .A2(_4358_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8338_ (.A1(_3502_),
    .A2(_3538_),
    .B(_3539_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8339_ (.A1(_0321_),
    .A2(_0326_),
    .B(_0347_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8340_ (.A1(_1404_),
    .A2(_0327_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8341_ (.A1(_3541_),
    .A2(_3542_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8342_ (.I(_4060_),
    .Z(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8343_ (.A1(_3540_),
    .A2(_3543_),
    .B(_3544_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8344_ (.A1(_3540_),
    .A2(_3543_),
    .B(_3545_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8345_ (.A1(_1404_),
    .A2(_3544_),
    .B(_3507_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8346_ (.A1(_1502_),
    .A2(_4374_),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8347_ (.A1(_3510_),
    .A2(_3511_),
    .B(_3548_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8348_ (.A1(_1403_),
    .A2(_0331_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8349_ (.A1(_3549_),
    .A2(_3550_),
    .B(_4097_),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8350_ (.A1(_3549_),
    .A2(_3550_),
    .B(_3551_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8351_ (.A1(_1404_),
    .A2(_3509_),
    .B(_3552_),
    .C(_2625_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8352_ (.A1(_3546_),
    .A2(_3547_),
    .B(_3553_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8353_ (.A1(_3472_),
    .A2(_3554_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8354_ (.A1(_3534_),
    .A2(_3536_),
    .B1(_3527_),
    .B2(_3537_),
    .C(_3555_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8355_ (.A1(_1473_),
    .A2(_3532_),
    .B1(_3556_),
    .B2(_3294_),
    .ZN(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8356_ (.A1(_1359_),
    .A2(_2490_),
    .B(_2485_),
    .ZN(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8357_ (.A1(_1623_),
    .A2(_3558_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8358_ (.A1(_3461_),
    .A2(_3557_),
    .B(_3559_),
    .C(_3485_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8359_ (.A1(net30),
    .A2(_3460_),
    .B(_3560_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8360_ (.A1(_3338_),
    .A2(_3561_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8361_ (.I(net31),
    .ZN(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8362_ (.A1(net30),
    .A2(net53),
    .A3(net28),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8363_ (.A1(_3562_),
    .A2(_3563_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8364_ (.I(_3465_),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8365_ (.A1(_0347_),
    .A2(_0321_),
    .A3(_0326_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8366_ (.A1(_3540_),
    .A2(_3541_),
    .B(_3566_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8367_ (.A1(_1484_),
    .A2(_0458_),
    .A3(_3567_),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8368_ (.A1(_3565_),
    .A2(_3568_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8369_ (.A1(_1406_),
    .A2(_3565_),
    .B(_3464_),
    .C(_3569_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8370_ (.I(_4097_),
    .Z(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8371_ (.I(_3571_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8372_ (.A1(_0348_),
    .A2(_0330_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8373_ (.A1(_0348_),
    .A2(_0330_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8374_ (.A1(_3549_),
    .A2(_3573_),
    .B(_3574_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8375_ (.A1(_1484_),
    .A2(_0452_),
    .A3(_3575_),
    .Z(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8376_ (.A1(_3571_),
    .A2(_3576_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8377_ (.A1(_1407_),
    .A2(_3572_),
    .B(_3577_),
    .C(_2622_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8378_ (.I(_2404_),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8379_ (.A1(_3570_),
    .A2(_3578_),
    .B(_3579_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8380_ (.A1(_3537_),
    .A2(_3564_),
    .B(_3580_),
    .C(_2629_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8381_ (.A1(_1621_),
    .A2(_1402_),
    .B(_3534_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8382_ (.A1(_2846_),
    .A2(_3582_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8383_ (.A1(_3500_),
    .A2(_3583_),
    .B(_3519_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8384_ (.A1(_2788_),
    .A2(_2849_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8385_ (.A1(_2897_),
    .A2(_3564_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8386_ (.A1(_2852_),
    .A2(_3586_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8387_ (.A1(_1256_),
    .A2(_2701_),
    .A3(_3587_),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8388_ (.A1(_1631_),
    .A2(_2548_),
    .A3(_2569_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8389_ (.A1(_1568_),
    .A2(_3588_),
    .A3(_3589_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8390_ (.A1(_1631_),
    .A2(_2586_),
    .B1(_3585_),
    .B2(_3590_),
    .ZN(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8391_ (.A1(_3581_),
    .A2(_3584_),
    .B(_3591_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8392_ (.A1(_1729_),
    .A2(_3490_),
    .B1(_3592_),
    .B2(_2572_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8393_ (.A1(net31),
    .A2(_3523_),
    .B(_3191_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8394_ (.A1(_3489_),
    .A2(_3593_),
    .B(_3594_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8395_ (.I(_2532_),
    .Z(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8396_ (.I(_2405_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8397_ (.A1(_3562_),
    .A2(_3563_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8398_ (.A1(net32),
    .A2(_3597_),
    .Z(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8399_ (.A1(_2845_),
    .A2(_3582_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8400_ (.A1(_2844_),
    .A2(_3599_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8401_ (.A1(_2887_),
    .A2(_3600_),
    .Z(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8402_ (.I(_2559_),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8403_ (.I(_3544_),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8404_ (.A1(_0430_),
    .A2(_0457_),
    .ZN(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _8405_ (.A1(_2899_),
    .A2(_0457_),
    .B1(_3540_),
    .B2(_3541_),
    .C(_3566_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8406_ (.A1(_3604_),
    .A2(_3605_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8407_ (.A1(_1409_),
    .A2(_0516_),
    .A3(_3606_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8408_ (.A1(_3603_),
    .A2(_3607_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8409_ (.A1(_1411_),
    .A2(_3603_),
    .B(_3507_),
    .C(_3608_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8410_ (.A1(_2899_),
    .A2(_0451_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _8411_ (.A1(_2899_),
    .A2(_0451_),
    .B1(_3549_),
    .B2(_3573_),
    .C(_3574_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8412_ (.A1(_3610_),
    .A2(_3611_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8413_ (.A1(_1409_),
    .A2(_0553_),
    .A3(_3612_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8414_ (.A1(_3509_),
    .A2(_3613_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8415_ (.A1(_1411_),
    .A2(_3509_),
    .B(_3614_),
    .C(_2626_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8416_ (.A1(_3609_),
    .A2(_3615_),
    .B(_3515_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8417_ (.A1(_3596_),
    .A2(_3598_),
    .B1(_3601_),
    .B2(_3602_),
    .C(_3616_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8418_ (.A1(_2851_),
    .A2(_3598_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8419_ (.A1(_2910_),
    .A2(_3618_),
    .B(_3492_),
    .ZN(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8420_ (.A1(_2884_),
    .A2(_2890_),
    .B(_3619_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8421_ (.A1(_1689_),
    .A2(_3525_),
    .B1(_3620_),
    .B2(_2473_),
    .C(_2687_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8422_ (.A1(_1639_),
    .A2(_3558_),
    .B(_3621_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8423_ (.A1(_2459_),
    .A2(_3617_),
    .B(_3622_),
    .C(_3485_),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8424_ (.A1(net32),
    .A2(_3460_),
    .B(_3623_),
    .ZN(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8425_ (.A1(_3595_),
    .A2(_3624_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8426_ (.I(_3488_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8427_ (.I(_2580_),
    .Z(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8428_ (.A1(_2887_),
    .A2(_3600_),
    .Z(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8429_ (.A1(_2933_),
    .A2(_3627_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8430_ (.A1(_2932_),
    .A2(_3628_),
    .Z(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8431_ (.A1(net32),
    .A2(_3597_),
    .Z(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8432_ (.A1(net52),
    .A2(_3630_),
    .Z(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8433_ (.A1(_0538_),
    .A2(_0515_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8434_ (.A1(_0539_),
    .A2(_0515_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8435_ (.A1(_3604_),
    .A2(_3632_),
    .A3(_3605_),
    .B(_3633_),
    .ZN(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8436_ (.A1(_0605_),
    .A2(_0619_),
    .Z(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8437_ (.A1(_3634_),
    .A2(_3635_),
    .B(_4060_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8438_ (.A1(_3634_),
    .A2(_3635_),
    .B(_3636_),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8439_ (.A1(_1282_),
    .A2(_3565_),
    .B(_2287_),
    .C(_3637_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8440_ (.I(_0603_),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8441_ (.A1(_3639_),
    .A2(_0587_),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8442_ (.A1(_3639_),
    .A2(_0586_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8443_ (.A1(_0538_),
    .A2(_0552_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8444_ (.A1(_0539_),
    .A2(_0552_),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8445_ (.A1(_3610_),
    .A2(_3642_),
    .A3(_3611_),
    .B(_3643_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8446_ (.A1(_3640_),
    .A2(_3641_),
    .A3(_3644_),
    .ZN(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8447_ (.A1(_3640_),
    .A2(_3641_),
    .B(_3644_),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8448_ (.A1(_3571_),
    .A2(_3646_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8449_ (.A1(_1282_),
    .A2(_3571_),
    .B1(_3645_),
    .B2(_3647_),
    .C(_2255_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8450_ (.A1(_3638_),
    .A2(_3648_),
    .B(_3579_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8451_ (.A1(_3537_),
    .A2(_3631_),
    .B(_3649_),
    .C(_2580_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8452_ (.A1(_3626_),
    .A2(_3629_),
    .B(_3650_),
    .C(_3294_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8453_ (.A1(_2868_),
    .A2(_3631_),
    .ZN(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8454_ (.A1(_2949_),
    .A2(_3652_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8455_ (.I(_2668_),
    .Z(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8456_ (.A1(_1644_),
    .A2(_3480_),
    .B1(_3653_),
    .B2(_3654_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8457_ (.A1(_2791_),
    .A2(_2936_),
    .A3(_3655_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8458_ (.A1(_1645_),
    .A2(_3484_),
    .B1(_3651_),
    .B2(_3461_),
    .C(_3656_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8459_ (.A1(net33),
    .A2(_3488_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8460_ (.I(_1294_),
    .Z(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8461_ (.A1(_3625_),
    .A2(_3657_),
    .B(_3658_),
    .C(_3659_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8462_ (.A1(net52),
    .A2(_3630_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8463_ (.A1(net34),
    .A2(_3660_),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8464_ (.A1(_2804_),
    .A2(_3661_),
    .B(_2980_),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8465_ (.A1(_3040_),
    .A2(_2975_),
    .B1(_3493_),
    .B2(_3662_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8466_ (.I(_3663_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8467_ (.A1(_1650_),
    .A2(_3491_),
    .B1(_3664_),
    .B2(_3498_),
    .ZN(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8468_ (.A1(_3463_),
    .A2(_3661_),
    .B(_3517_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8469_ (.A1(_0725_),
    .A2(_0708_),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8470_ (.I(_3641_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8471_ (.A1(_3640_),
    .A2(_3644_),
    .B(_3668_),
    .ZN(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8472_ (.A1(_3667_),
    .A2(_3669_),
    .B(_3468_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8473_ (.A1(_3667_),
    .A2(_3669_),
    .B(_3670_),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8474_ (.A1(_1412_),
    .A2(_3572_),
    .B(_3671_),
    .C(_2622_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8475_ (.A1(_0725_),
    .A2(_0734_),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8476_ (.A1(_3639_),
    .A2(_0618_),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8477_ (.A1(_3639_),
    .A2(_0618_),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8478_ (.A1(_3634_),
    .A2(_3674_),
    .B(_3675_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8479_ (.A1(_3673_),
    .A2(_3676_),
    .Z(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8480_ (.A1(_0726_),
    .A2(_3544_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8481_ (.A1(_3603_),
    .A2(_3677_),
    .B(_3678_),
    .C(_2287_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8482_ (.A1(_3672_),
    .A2(_3679_),
    .B(_3579_),
    .ZN(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8483_ (.A1(_2932_),
    .A2(_3627_),
    .B(_2973_),
    .ZN(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8484_ (.A1(_2970_),
    .A2(_3681_),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8485_ (.A1(_3666_),
    .A2(_3680_),
    .B1(_3682_),
    .B2(_3500_),
    .C(_3473_),
    .ZN(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8486_ (.A1(_1360_),
    .A2(_3665_),
    .B(_3683_),
    .ZN(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8487_ (.A1(_1696_),
    .A2(_3490_),
    .B1(_3684_),
    .B2(_2572_),
    .ZN(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8488_ (.A1(net34),
    .A2(_3523_),
    .B(_3191_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8489_ (.A1(_3489_),
    .A2(_3685_),
    .B(_3686_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8490_ (.A1(_1372_),
    .A2(_0709_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8491_ (.A1(_3667_),
    .A2(_3669_),
    .B(_3687_),
    .ZN(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8492_ (.A1(_1519_),
    .A2(_0781_),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8493_ (.A1(_3688_),
    .A2(_3689_),
    .B(_3572_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8494_ (.A1(_3688_),
    .A2(_3689_),
    .B(_3690_),
    .ZN(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8495_ (.A1(_1393_),
    .A2(_3572_),
    .B(_2482_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8496_ (.A1(_1491_),
    .A2(_0735_),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8497_ (.A1(_3673_),
    .A2(_3676_),
    .B(_3693_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8498_ (.A1(_1519_),
    .A2(_0797_),
    .A3(_3694_),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8499_ (.A1(_3603_),
    .A2(_3695_),
    .ZN(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8500_ (.A1(_1393_),
    .A2(_3565_),
    .B(_3464_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8501_ (.A1(_3691_),
    .A2(_3692_),
    .B1(_3696_),
    .B2(_3697_),
    .ZN(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8502_ (.A1(net34),
    .A2(net52),
    .A3(_3630_),
    .ZN(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8503_ (.A1(net35),
    .A2(_3699_),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8504_ (.A1(_3596_),
    .A2(_3700_),
    .ZN(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8505_ (.A1(_3515_),
    .A2(_3698_),
    .B(_3701_),
    .C(_3626_),
    .ZN(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8506_ (.A1(_2970_),
    .A2(_3681_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8507_ (.A1(_3021_),
    .A2(_3703_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8508_ (.A1(_3020_),
    .A2(_3704_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8509_ (.A1(_3602_),
    .A2(_3705_),
    .B(_2459_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8510_ (.A1(_3702_),
    .A2(_3706_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8511_ (.A1(_2558_),
    .A2(_2862_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8512_ (.A1(_3326_),
    .A2(_3700_),
    .B(_3708_),
    .ZN(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8513_ (.A1(_1656_),
    .A2(_3491_),
    .B1(_3709_),
    .B2(_3654_),
    .C(_3042_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8514_ (.A1(_2732_),
    .A2(_3710_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8515_ (.A1(_1657_),
    .A2(_3484_),
    .B(_3707_),
    .C(_3711_),
    .ZN(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8516_ (.I(_3459_),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8517_ (.I(_2338_),
    .Z(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8518_ (.A1(net35),
    .A2(_3713_),
    .B(_3714_),
    .ZN(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8519_ (.A1(_3489_),
    .A2(_3712_),
    .B(_3715_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8520_ (.I(net36),
    .Z(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8521_ (.I(net35),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8522_ (.A1(_3717_),
    .A2(_3699_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8523_ (.A1(_3716_),
    .A2(_3718_),
    .ZN(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8524_ (.A1(_2252_),
    .A2(_3326_),
    .ZN(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8525_ (.A1(_3326_),
    .A2(_3719_),
    .B(_3493_),
    .C(_3720_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8526_ (.A1(_2470_),
    .A2(_3058_),
    .B(_3721_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8527_ (.A1(_3051_),
    .A2(_3491_),
    .B1(_3722_),
    .B2(_3498_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8528_ (.A1(_0783_),
    .A2(_0780_),
    .ZN(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8529_ (.A1(_3667_),
    .A2(_3669_),
    .B(_3724_),
    .C(_3687_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8530_ (.A1(_1488_),
    .A2(_0780_),
    .ZN(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8531_ (.A1(_4097_),
    .A2(_3726_),
    .ZN(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8532_ (.A1(_3725_),
    .A2(_3727_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8533_ (.A1(_2252_),
    .A2(_3728_),
    .Z(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8534_ (.A1(_0783_),
    .A2(_0796_),
    .ZN(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8535_ (.A1(_3673_),
    .A2(_3676_),
    .B(_3730_),
    .C(_3693_),
    .ZN(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8536_ (.A1(_1488_),
    .A2(_0796_),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8537_ (.A1(_4365_),
    .A2(_3732_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8538_ (.A1(_3731_),
    .A2(_3733_),
    .ZN(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8539_ (.A1(_2252_),
    .A2(_3734_),
    .Z(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8540_ (.A1(_3340_),
    .A2(_3729_),
    .B1(_3735_),
    .B2(_3507_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8541_ (.A1(_3596_),
    .A2(_3719_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8542_ (.A1(_3515_),
    .A2(_3736_),
    .B(_3737_),
    .C(_3626_),
    .ZN(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8543_ (.A1(_3055_),
    .A2(_3681_),
    .B(_3056_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8544_ (.A1(_3054_),
    .A2(_3739_),
    .Z(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8545_ (.A1(_3054_),
    .A2(_3739_),
    .B(_2629_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8546_ (.A1(_3740_),
    .A2(_3741_),
    .B(_2458_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8547_ (.A1(_3051_),
    .A2(_3558_),
    .B1(_3738_),
    .B2(_3742_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8548_ (.A1(_2831_),
    .A2(_3723_),
    .B(_3743_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8549_ (.A1(_3716_),
    .A2(_3713_),
    .B(_3714_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8550_ (.A1(_3625_),
    .A2(_3744_),
    .B(_3745_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8551_ (.A1(_3089_),
    .A2(_3740_),
    .ZN(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8552_ (.A1(_3088_),
    .A2(_3746_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8553_ (.A1(_3062_),
    .A2(_3731_),
    .A3(_3733_),
    .ZN(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8554_ (.A1(_2296_),
    .A2(_3748_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8555_ (.A1(_3062_),
    .A2(_3725_),
    .A3(_3727_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8556_ (.A1(_3097_),
    .A2(_3750_),
    .ZN(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8557_ (.A1(_3464_),
    .A2(_3749_),
    .B1(_3751_),
    .B2(_2256_),
    .ZN(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8558_ (.A1(_3716_),
    .A2(_3718_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8559_ (.A1(net51),
    .A2(_3753_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8560_ (.A1(_3579_),
    .A2(_3752_),
    .B1(_3754_),
    .B2(_3463_),
    .C(_3517_),
    .ZN(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8561_ (.A1(_3602_),
    .A2(_3747_),
    .B(_3755_),
    .C(_2459_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8562_ (.A1(_2862_),
    .A2(_3754_),
    .B(_3098_),
    .ZN(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8563_ (.A1(_1106_),
    .A2(_3525_),
    .B1(_3757_),
    .B2(_3654_),
    .C(_2437_),
    .ZN(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8564_ (.A1(_3093_),
    .A2(_3758_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8565_ (.A1(_1106_),
    .A2(_3484_),
    .B(_3759_),
    .ZN(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8566_ (.A1(_3756_),
    .A2(_3760_),
    .B(_3488_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8567_ (.A1(net51),
    .A2(_3460_),
    .B(_3761_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8568_ (.A1(_3595_),
    .A2(_3762_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8569_ (.A1(_3472_),
    .A2(_2286_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8570_ (.A1(_3063_),
    .A2(_2296_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8571_ (.A1(_3725_),
    .A2(_3727_),
    .B(_4092_),
    .ZN(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8572_ (.A1(_3731_),
    .A2(_3733_),
    .B(_2561_),
    .ZN(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8573_ (.A1(_3764_),
    .A2(_3765_),
    .A3(_3766_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8574_ (.A1(_2298_),
    .A2(_3767_),
    .Z(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8575_ (.A1(net51),
    .A2(net36),
    .A3(_3718_),
    .ZN(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8576_ (.A1(net38),
    .A2(_3769_),
    .ZN(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8577_ (.A1(_3505_),
    .A2(_3770_),
    .Z(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8578_ (.A1(_3763_),
    .A2(_3768_),
    .B(_3771_),
    .C(_2629_),
    .ZN(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8579_ (.A1(_3088_),
    .A2(_3740_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8580_ (.A1(_3123_),
    .A2(_3773_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8581_ (.A1(_3120_),
    .A2(_3774_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8582_ (.A1(_3500_),
    .A2(_3775_),
    .B(_3519_),
    .ZN(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8583_ (.A1(_2546_),
    .A2(_3770_),
    .ZN(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8584_ (.A1(_3126_),
    .A2(_3777_),
    .ZN(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8585_ (.A1(_3040_),
    .A2(_3125_),
    .B1(_3493_),
    .B2(_3778_),
    .ZN(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8586_ (.I(_3779_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8587_ (.A1(_1114_),
    .A2(_3480_),
    .B1(_3780_),
    .B2(_3498_),
    .ZN(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8588_ (.A1(_3772_),
    .A2(_3776_),
    .B1(_3781_),
    .B2(_1360_),
    .ZN(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8589_ (.A1(_1114_),
    .A2(_3490_),
    .B1(_3782_),
    .B2(_3461_),
    .ZN(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8590_ (.A1(net38),
    .A2(_3713_),
    .B(_3714_),
    .ZN(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8591_ (.A1(_3625_),
    .A2(_3783_),
    .B(_3784_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8592_ (.A1(_2301_),
    .A2(_3144_),
    .A3(_3765_),
    .A4(_3766_),
    .Z(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8593_ (.A1(_3144_),
    .A2(_3766_),
    .B(_2301_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8594_ (.A1(_3785_),
    .A2(_3786_),
    .B(_3506_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8595_ (.A1(_3144_),
    .A2(_3728_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8596_ (.A1(_3143_),
    .A2(_2482_),
    .A3(_3788_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8597_ (.A1(_3787_),
    .A2(_3789_),
    .B(_3472_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8598_ (.A1(net38),
    .A2(net51),
    .A3(_3716_),
    .A4(_3718_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8599_ (.A1(net39),
    .A2(_3791_),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8600_ (.A1(_3596_),
    .A2(_3792_),
    .B(_2620_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8601_ (.A1(_3120_),
    .A2(_3774_),
    .B(_3148_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8602_ (.A1(_3147_),
    .A2(_3794_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8603_ (.A1(_3790_),
    .A2(_3793_),
    .B1(_3795_),
    .B2(_3602_),
    .C(_2458_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8604_ (.A1(_2892_),
    .A2(_3150_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8605_ (.A1(_2862_),
    .A2(_3792_),
    .B(_3151_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8606_ (.A1(_1122_),
    .A2(_3525_),
    .B1(_3798_),
    .B2(_2668_),
    .C(_2437_),
    .ZN(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8607_ (.A1(_3797_),
    .A2(_3799_),
    .ZN(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8608_ (.A1(_1122_),
    .A2(_3483_),
    .B(_3800_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8609_ (.A1(_3796_),
    .A2(_3801_),
    .B(_3485_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8610_ (.A1(net39),
    .A2(_3523_),
    .B(_3802_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8611_ (.A1(_3595_),
    .A2(_3803_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8612_ (.A1(_2306_),
    .A2(_3785_),
    .Z(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8613_ (.I(net39),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8614_ (.A1(_3805_),
    .A2(_3791_),
    .ZN(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8615_ (.A1(net40),
    .A2(_3806_),
    .Z(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8616_ (.A1(_3537_),
    .A2(_3804_),
    .B1(_3807_),
    .B2(_3763_),
    .C(_2620_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8617_ (.A1(_3169_),
    .A2(_3773_),
    .B(_3171_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8618_ (.A1(_3173_),
    .A2(_3809_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8619_ (.A1(_3626_),
    .A2(_3810_),
    .ZN(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8620_ (.A1(_2898_),
    .A2(_3807_),
    .ZN(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8621_ (.A1(_3180_),
    .A2(_3812_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8622_ (.A1(_1130_),
    .A2(_3480_),
    .B1(_3813_),
    .B2(_3654_),
    .C(_3175_),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8623_ (.A1(_3519_),
    .A2(_3808_),
    .A3(_3811_),
    .B1(_3814_),
    .B2(_2481_),
    .ZN(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8624_ (.A1(_1130_),
    .A2(_3558_),
    .B1(_3815_),
    .B2(_2485_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8625_ (.A1(net40),
    .A2(_3713_),
    .B(_3714_),
    .ZN(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8626_ (.A1(_3625_),
    .A2(_3816_),
    .B(_3817_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8627_ (.A1(_0967_),
    .A2(_1145_),
    .ZN(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8628_ (.I(_3818_),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8629_ (.I(_3819_),
    .Z(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8630_ (.I(_3819_),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8631_ (.A1(\as2650.stack[4][8] ),
    .A2(_3821_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8632_ (.A1(_1190_),
    .A2(_3820_),
    .B(_3822_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8633_ (.I(_3818_),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8634_ (.A1(\as2650.stack[4][9] ),
    .A2(_3823_),
    .ZN(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8635_ (.A1(_1200_),
    .A2(_3820_),
    .B(_3824_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8636_ (.A1(\as2650.stack[4][10] ),
    .A2(_3823_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8637_ (.A1(_1203_),
    .A2(_3820_),
    .B(_3825_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8638_ (.A1(\as2650.stack[4][11] ),
    .A2(_3823_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8639_ (.A1(_1205_),
    .A2(_3820_),
    .B(_3826_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8640_ (.A1(\as2650.stack[4][12] ),
    .A2(_3823_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8641_ (.A1(_1207_),
    .A2(_3821_),
    .B(_3827_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8642_ (.A1(\as2650.stack[4][13] ),
    .A2(_3819_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8643_ (.A1(_1209_),
    .A2(_3821_),
    .B(_3828_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8644_ (.A1(\as2650.stack[4][14] ),
    .A2(_3819_),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8645_ (.A1(_1211_),
    .A2(_3821_),
    .B(_3829_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8646_ (.I(net41),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8647_ (.A1(_2253_),
    .A2(_2317_),
    .A3(_2411_),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8648_ (.A1(_0940_),
    .A2(_2571_),
    .A3(_2673_),
    .ZN(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8649_ (.A1(_1214_),
    .A2(_2319_),
    .ZN(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8650_ (.A1(_4195_),
    .A2(_2350_),
    .B(_3234_),
    .C(_3833_),
    .ZN(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8651_ (.A1(_3223_),
    .A2(_3831_),
    .A3(_3832_),
    .A4(_3834_),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8652_ (.I(_3835_),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8653_ (.I(_0864_),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8654_ (.I(_3837_),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8655_ (.I(_3835_),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8656_ (.I(_3837_),
    .Z(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8657_ (.A1(_1589_),
    .A2(_3840_),
    .ZN(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8658_ (.A1(_3838_),
    .A2(_3262_),
    .B(_3839_),
    .C(_3841_),
    .ZN(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8659_ (.A1(_3830_),
    .A2(_3836_),
    .B(_3842_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8660_ (.I(_3837_),
    .Z(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8661_ (.A1(_1610_),
    .A2(_3843_),
    .ZN(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8662_ (.A1(_3838_),
    .A2(_3258_),
    .B(_3844_),
    .ZN(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8663_ (.I(_3835_),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8664_ (.A1(net42),
    .A2(_3846_),
    .ZN(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8665_ (.A1(_3836_),
    .A2(_3845_),
    .B(_3847_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8666_ (.A1(_1619_),
    .A2(_3843_),
    .ZN(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8667_ (.A1(_3838_),
    .A2(_2014_),
    .B(_3848_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8668_ (.A1(net43),
    .A2(_3846_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8669_ (.A1(_3836_),
    .A2(_3849_),
    .B(_3850_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8670_ (.I(_3835_),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8671_ (.I(_3837_),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8672_ (.A1(_1628_),
    .A2(_3843_),
    .ZN(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8673_ (.A1(_3852_),
    .A2(_1388_),
    .B(_3853_),
    .ZN(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8674_ (.A1(net44),
    .A2(_3846_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8675_ (.A1(_3851_),
    .A2(_3854_),
    .B(_3855_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8676_ (.A1(_1635_),
    .A2(_3843_),
    .ZN(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8677_ (.A1(_3852_),
    .A2(_0591_),
    .B(_3856_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8678_ (.A1(net45),
    .A2(_3846_),
    .ZN(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8679_ (.A1(_3851_),
    .A2(_3857_),
    .B(_3858_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8680_ (.I(net19),
    .ZN(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8681_ (.A1(_0590_),
    .A2(_3840_),
    .ZN(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8682_ (.A1(_3838_),
    .A2(_0646_),
    .B(_3839_),
    .C(_3860_),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8683_ (.A1(_3859_),
    .A2(_3836_),
    .B(_3861_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8684_ (.A1(_0713_),
    .A2(_3840_),
    .ZN(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8685_ (.A1(_3852_),
    .A2(_0681_),
    .B(_3862_),
    .ZN(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8686_ (.A1(net20),
    .A2(_3839_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8687_ (.A1(_3851_),
    .A2(_3863_),
    .B(_3864_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8688_ (.A1(_1040_),
    .A2(_3840_),
    .ZN(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8689_ (.A1(_3852_),
    .A2(_0717_),
    .B(_3865_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8690_ (.A1(net21),
    .A2(_3839_),
    .ZN(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8691_ (.A1(_3851_),
    .A2(_3866_),
    .B(_3867_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8692_ (.A1(_2303_),
    .A2(_1573_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8693_ (.A1(_2431_),
    .A2(_1576_),
    .B(_3868_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8694_ (.I(_2267_),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8695_ (.A1(_2307_),
    .A2(_1573_),
    .ZN(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8696_ (.A1(_3869_),
    .A2(_1576_),
    .B(_3870_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8697_ (.A1(_2354_),
    .A2(_1227_),
    .A3(_1245_),
    .A4(_2314_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8698_ (.A1(_2658_),
    .A2(_1461_),
    .A3(_2400_),
    .A4(_3871_),
    .ZN(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8699_ (.A1(_1432_),
    .A2(_3872_),
    .ZN(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8700_ (.A1(_0403_),
    .A2(_1846_),
    .ZN(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8701_ (.A1(_1464_),
    .A2(_1544_),
    .ZN(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8702_ (.A1(_1445_),
    .A2(_2317_),
    .A3(_3874_),
    .A4(_3875_),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8703_ (.A1(_0939_),
    .A2(_2324_),
    .A3(_3876_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8704_ (.A1(_1457_),
    .A2(_1458_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8705_ (.A1(_4207_),
    .A2(_1859_),
    .B1(_1220_),
    .B2(_2280_),
    .C(_3878_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8706_ (.A1(_3873_),
    .A2(_3877_),
    .A3(_3879_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8707_ (.A1(_1283_),
    .A2(_2550_),
    .A3(_2677_),
    .ZN(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8708_ (.A1(_3880_),
    .A2(_3881_),
    .ZN(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8709_ (.A1(_1266_),
    .A2(_1280_),
    .ZN(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8710_ (.A1(_1528_),
    .A2(_2522_),
    .A3(_3883_),
    .ZN(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8711_ (.A1(_3344_),
    .A2(_3884_),
    .B(_3313_),
    .ZN(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8712_ (.A1(_3313_),
    .A2(_0681_),
    .B(_3885_),
    .ZN(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8713_ (.A1(_2481_),
    .A2(_0511_),
    .ZN(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8714_ (.A1(_3869_),
    .A2(_3886_),
    .B(_3882_),
    .C(_3887_),
    .ZN(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8715_ (.A1(\as2650.psl[5] ),
    .A2(_3882_),
    .B(_3888_),
    .ZN(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8716_ (.A1(_3595_),
    .A2(_3889_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8717_ (.A1(_0639_),
    .A2(_2096_),
    .ZN(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8718_ (.A1(_0407_),
    .A2(_0412_),
    .ZN(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8719_ (.A1(_0640_),
    .A2(_0355_),
    .ZN(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8720_ (.A1(_0387_),
    .A2(_2493_),
    .B(_3892_),
    .ZN(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8721_ (.A1(_0315_),
    .A2(_3893_),
    .ZN(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8722_ (.A1(_4325_),
    .A2(_4159_),
    .ZN(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8723_ (.A1(_0486_),
    .A2(_4184_),
    .B(_3895_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8724_ (.A1(_4329_),
    .A2(_4353_),
    .B(_4169_),
    .C(_3896_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8725_ (.A1(_4329_),
    .A2(_4354_),
    .ZN(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8726_ (.A1(_0315_),
    .A2(_3893_),
    .B(_3897_),
    .C(_3898_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8727_ (.A1(_3891_),
    .A2(_3894_),
    .A3(_3899_),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8728_ (.A1(_0407_),
    .A2(_0413_),
    .B1(_0628_),
    .B2(_0510_),
    .C(_3900_),
    .ZN(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8729_ (.A1(_0488_),
    .A2(_0509_),
    .B1(_0639_),
    .B2(_2096_),
    .C(_3901_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8730_ (.A1(_0692_),
    .A2(_0701_),
    .ZN(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8731_ (.A1(_3890_),
    .A2(_3902_),
    .B(_3903_),
    .ZN(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8732_ (.A1(_2493_),
    .A2(_1340_),
    .ZN(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8733_ (.A1(\as2650.holding_reg[7] ),
    .A2(_2493_),
    .B(_3905_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8734_ (.A1(_0692_),
    .A2(_0701_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8735_ (.A1(_1311_),
    .A2(_3906_),
    .B(_3907_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8736_ (.A1(_1311_),
    .A2(_3906_),
    .ZN(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8737_ (.A1(_3904_),
    .A2(_3908_),
    .B(_3909_),
    .C(_3869_),
    .ZN(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8738_ (.I(_1266_),
    .Z(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8739_ (.A1(_3911_),
    .A2(_2488_),
    .B(_3303_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8740_ (.A1(_3303_),
    .A2(_0717_),
    .B1(_2492_),
    .B2(_3912_),
    .C(_3313_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8741_ (.A1(_1383_),
    .A2(_3262_),
    .B(_1362_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8742_ (.A1(_1399_),
    .A2(_2550_),
    .A3(_2677_),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8743_ (.A1(_3880_),
    .A2(_3915_),
    .ZN(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8744_ (.A1(_3913_),
    .A2(_3914_),
    .B(_3916_),
    .ZN(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8745_ (.I(_3917_),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8746_ (.A1(\as2650.carry ),
    .A2(_3916_),
    .B(_2534_),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8747_ (.A1(_3910_),
    .A2(_3918_),
    .B(_3919_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8748_ (.I(_2421_),
    .Z(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8749_ (.A1(_2299_),
    .A2(_3920_),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8750_ (.A1(_1228_),
    .A2(_1250_),
    .B(_2335_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8751_ (.I(_2669_),
    .ZN(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8752_ (.A1(_2664_),
    .A2(_3923_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8753_ (.A1(_1237_),
    .A2(_2676_),
    .B(_1424_),
    .ZN(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8754_ (.A1(_2542_),
    .A2(_2325_),
    .A3(_2598_),
    .ZN(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8755_ (.A1(_2257_),
    .A2(_3926_),
    .ZN(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8756_ (.A1(_4314_),
    .A2(_3251_),
    .ZN(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8757_ (.A1(_4308_),
    .A2(_3928_),
    .B(_2706_),
    .C(_2646_),
    .ZN(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8758_ (.A1(_2530_),
    .A2(_3282_),
    .ZN(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8759_ (.A1(_1273_),
    .A2(_1068_),
    .B(_2467_),
    .C(_3930_),
    .ZN(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8760_ (.A1(_1500_),
    .A2(_1259_),
    .B(_2883_),
    .ZN(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8761_ (.A1(_1265_),
    .A2(_1464_),
    .A3(_2480_),
    .A4(_3932_),
    .ZN(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8762_ (.A1(_3927_),
    .A2(_3929_),
    .A3(_3931_),
    .A4(_3933_),
    .ZN(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _8763_ (.A1(_3922_),
    .A2(_3924_),
    .A3(_3925_),
    .A4(_3934_),
    .Z(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8764_ (.A1(_3921_),
    .A2(_3935_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8765_ (.I(_2603_),
    .Z(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8766_ (.A1(_1713_),
    .A2(_1048_),
    .Z(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8767_ (.A1(_0334_),
    .A2(_1092_),
    .ZN(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8768_ (.I(_1261_),
    .Z(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8769_ (.A1(_3940_),
    .A2(_3938_),
    .ZN(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8770_ (.A1(_1355_),
    .A2(_3253_),
    .A3(_3939_),
    .A4(_3941_),
    .ZN(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8771_ (.A1(_1575_),
    .A2(_1288_),
    .B(_1336_),
    .ZN(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8772_ (.A1(_3942_),
    .A2(_3943_),
    .ZN(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8773_ (.A1(_0965_),
    .A2(_1279_),
    .ZN(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8774_ (.A1(_1279_),
    .A2(_3944_),
    .B1(_3945_),
    .B2(_0957_),
    .C(_3937_),
    .ZN(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8775_ (.A1(_3937_),
    .A2(_3938_),
    .B(_3946_),
    .ZN(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8776_ (.A1(_1747_),
    .A2(_3936_),
    .B(_2534_),
    .ZN(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8777_ (.A1(_3936_),
    .A2(_3947_),
    .B(_3948_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8778_ (.A1(_1572_),
    .A2(_3920_),
    .ZN(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8779_ (.A1(_3935_),
    .A2(_3949_),
    .ZN(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8780_ (.A1(_0892_),
    .A2(_0899_),
    .ZN(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8781_ (.A1(_1355_),
    .A2(_2657_),
    .ZN(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8782_ (.A1(_3951_),
    .A2(_1261_),
    .ZN(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8783_ (.A1(_1610_),
    .A2(_3940_),
    .B(_3953_),
    .ZN(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8784_ (.A1(_2428_),
    .A2(_0881_),
    .A3(_3954_),
    .ZN(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8785_ (.A1(_2505_),
    .A2(_3952_),
    .A3(_3955_),
    .B(_1279_),
    .ZN(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8786_ (.A1(_3951_),
    .A2(_3945_),
    .B(_3937_),
    .ZN(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8787_ (.A1(_3937_),
    .A2(_3951_),
    .B1(_3956_),
    .B2(_3957_),
    .ZN(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8788_ (.A1(_0902_),
    .A2(_3950_),
    .ZN(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8789_ (.A1(_3950_),
    .A2(_3958_),
    .B(_3959_),
    .C(_3659_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8790_ (.A1(_1559_),
    .A2(_3920_),
    .ZN(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8791_ (.A1(_3935_),
    .A2(_3960_),
    .ZN(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8792_ (.A1(_0947_),
    .A2(_3940_),
    .A3(_2488_),
    .B1(_2491_),
    .B2(_1288_),
    .ZN(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8793_ (.A1(_0881_),
    .A2(_3940_),
    .A3(_2996_),
    .ZN(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8794_ (.A1(_0905_),
    .A2(_3963_),
    .ZN(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8795_ (.A1(_2832_),
    .A2(_3962_),
    .B1(_3964_),
    .B2(_3920_),
    .ZN(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8796_ (.A1(_0905_),
    .A2(_3961_),
    .ZN(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8797_ (.A1(_3961_),
    .A2(_3965_),
    .B(_3966_),
    .C(_3659_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8798_ (.A1(_1405_),
    .A2(_2677_),
    .ZN(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8799_ (.A1(_1859_),
    .A2(_1220_),
    .A3(_3967_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8800_ (.A1(_3873_),
    .A2(_3877_),
    .A3(_3968_),
    .ZN(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8801_ (.A1(_3911_),
    .A2(_2510_),
    .B(_2509_),
    .ZN(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8802_ (.A1(_1474_),
    .A2(_3970_),
    .B(_3969_),
    .ZN(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8803_ (.A1(_1475_),
    .A2(_3906_),
    .Z(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8804_ (.A1(_3869_),
    .A2(_0803_),
    .A3(_3972_),
    .ZN(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8805_ (.A1(_1506_),
    .A2(_3969_),
    .B1(_3971_),
    .B2(_3973_),
    .C(_2639_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8806_ (.A1(_1258_),
    .A2(_1416_),
    .ZN(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _8807_ (.A1(_1553_),
    .A2(_1370_),
    .B(_2530_),
    .C(_2548_),
    .ZN(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8808_ (.A1(_1560_),
    .A2(_1500_),
    .ZN(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8809_ (.A1(_1258_),
    .A2(_1260_),
    .B(_1263_),
    .C(_3976_),
    .ZN(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8810_ (.A1(_1435_),
    .A2(_3974_),
    .A3(_3975_),
    .A4(_3977_),
    .ZN(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8811_ (.A1(_2307_),
    .A2(_2517_),
    .B(_3978_),
    .ZN(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8812_ (.A1(_2374_),
    .A2(_3976_),
    .ZN(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _8813_ (.A1(_1264_),
    .A2(_3975_),
    .A3(_3980_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8814_ (.A1(_2504_),
    .A2(_3911_),
    .B(_3974_),
    .C(_3981_),
    .ZN(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8815_ (.A1(_4286_),
    .A2(_3979_),
    .B1(_3982_),
    .B2(_2519_),
    .ZN(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8816_ (.A1(_2533_),
    .A2(_3983_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8817_ (.A1(_2303_),
    .A2(_2517_),
    .B(_3978_),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8818_ (.A1(_2515_),
    .A2(_3982_),
    .B1(_3984_),
    .B2(_4206_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8819_ (.A1(_2533_),
    .A2(_3985_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8820_ (.A1(_1572_),
    .A2(_2504_),
    .A3(_3911_),
    .ZN(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8821_ (.A1(_1777_),
    .A2(_2504_),
    .B(_3986_),
    .ZN(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8822_ (.A1(_2506_),
    .A2(_3978_),
    .B(\as2650.psl[1] ),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8823_ (.A1(_3978_),
    .A2(_3987_),
    .B(_3988_),
    .C(_3659_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8824_ (.A1(_1261_),
    .A2(_1221_),
    .A3(_3249_),
    .ZN(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8825_ (.A1(_1542_),
    .A2(_4311_),
    .A3(_3975_),
    .ZN(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8826_ (.A1(_2490_),
    .A2(_3989_),
    .B(_3990_),
    .ZN(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8827_ (.I(_3991_),
    .Z(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8828_ (.A1(_1584_),
    .A2(_3952_),
    .B(_2524_),
    .ZN(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8829_ (.A1(_2525_),
    .A2(_3992_),
    .B(_1492_),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8830_ (.A1(_3992_),
    .A2(_3993_),
    .B(_3994_),
    .ZN(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8831_ (.A1(_2533_),
    .A2(_3995_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8832_ (.A1(_2518_),
    .A2(_3992_),
    .B(\as2650.psu[4] ),
    .ZN(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8833_ (.A1(_3952_),
    .A2(_3991_),
    .ZN(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8834_ (.A1(_2519_),
    .A2(_3997_),
    .ZN(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8835_ (.A1(_3996_),
    .A2(_3998_),
    .B(_3049_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8836_ (.A1(_2514_),
    .A2(_3992_),
    .B(\as2650.psu[3] ),
    .ZN(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8837_ (.A1(_2515_),
    .A2(_3997_),
    .ZN(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8838_ (.A1(_3999_),
    .A2(_4000_),
    .B(_3049_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8839_ (.D(_0000_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8840_ (.D(_0001_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8841_ (.D(_0002_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8842_ (.D(_0003_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8843_ (.D(_0004_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8844_ (.D(_0005_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8845_ (.D(_0006_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8846_ (.D(_0007_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8847_ (.D(_0008_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8848_ (.D(_0009_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8849_ (.D(_0010_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8850_ (.D(_0011_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8851_ (.D(_0012_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8852_ (.D(_0013_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8853_ (.D(_0014_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8854_ (.D(_0015_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8855_ (.D(_0016_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8856_ (.D(_0017_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8857_ (.D(_0018_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8858_ (.D(_0019_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8859_ (.D(_0020_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8860_ (.D(_0021_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8861_ (.D(_0022_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8862_ (.D(_0023_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8863_ (.D(_0024_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8864_ (.D(_0025_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8865_ (.D(_0026_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8866_ (.D(_0027_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8867_ (.D(_0028_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8868_ (.D(_0029_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8869_ (.D(_0030_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8870_ (.D(_0031_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8871_ (.D(_0032_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8872_ (.D(_0033_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8873_ (.D(_0034_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8874_ (.D(_0035_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8875_ (.D(_0036_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8876_ (.D(_0037_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8877_ (.D(_0038_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8878_ (.D(_0039_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8879_ (.D(_0040_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8880_ (.D(_0041_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8881_ (.D(_0042_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8882_ (.D(_0043_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8883_ (.D(_0044_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8884_ (.D(_0045_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8885_ (.D(_0046_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8886_ (.D(_0047_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8887_ (.D(_0048_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8888_ (.D(_0049_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8889_ (.D(_0050_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8890_ (.D(_0051_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8891_ (.D(_0052_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8892_ (.D(_0053_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8893_ (.D(_0054_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8894_ (.D(_0055_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8895_ (.D(_0056_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8896_ (.D(_0057_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8897_ (.D(_0058_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8898_ (.D(_0059_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8899_ (.D(_0060_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8900_ (.D(_0061_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8901_ (.D(_0062_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8902_ (.D(_0063_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8903_ (.D(_0064_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8904_ (.D(_0065_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8905_ (.D(_0066_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8906_ (.D(_0067_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8907_ (.D(_0068_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8908_ (.D(_0069_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8909_ (.D(_0070_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8910_ (.D(_0071_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8911_ (.D(_0072_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8912_ (.D(_0073_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8913_ (.D(_0074_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8914_ (.D(_0075_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8915_ (.D(_0076_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8916_ (.D(_0077_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8917_ (.D(_0078_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8918_ (.D(_0079_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8919_ (.D(_0080_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8920_ (.D(_0081_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8921_ (.D(_0082_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8922_ (.D(_0083_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8923_ (.D(_0084_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8924_ (.D(_0085_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8925_ (.D(_0086_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8926_ (.D(_0087_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8927_ (.D(_0088_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8928_ (.D(_0089_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8929_ (.D(_0090_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8930_ (.D(_0091_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8931_ (.D(_0092_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8932_ (.D(_0093_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8933_ (.D(_0094_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8934_ (.D(_0095_),
    .CLK(clknet_opt_2_0_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8935_ (.D(_0096_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8936_ (.D(_0097_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8937_ (.D(_0098_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8938_ (.D(_0099_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8939_ (.D(_0100_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8940_ (.D(_0101_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8941_ (.D(_0102_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8942_ (.D(_0103_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8943_ (.D(_0104_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8944_ (.D(_0105_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8945_ (.D(_0106_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8946_ (.D(_0107_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8947_ (.D(_0108_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8948_ (.D(_0109_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8949_ (.D(_0110_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8950_ (.D(_0111_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8951_ (.D(_0112_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8952_ (.D(_0113_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8953_ (.D(_0114_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8954_ (.D(_0115_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8955_ (.D(_0116_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8956_ (.D(_0117_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8957_ (.D(_0118_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8958_ (.D(_0119_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8959_ (.D(_0120_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8960_ (.D(_0121_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8961_ (.D(_0122_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8962_ (.D(_0123_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8963_ (.D(_0124_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8964_ (.D(_0125_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8965_ (.D(_0126_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8966_ (.D(_0127_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8967_ (.D(_0128_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8968_ (.D(_0129_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8969_ (.D(_0130_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8970_ (.D(_0131_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8971_ (.D(_0132_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8972_ (.D(_0133_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8973_ (.D(_0134_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8974_ (.D(_0135_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8975_ (.D(_0136_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8976_ (.D(_0137_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8977_ (.D(_0138_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8978_ (.D(_0139_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8979_ (.D(_0140_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8980_ (.D(_0141_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8981_ (.D(_0142_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8982_ (.D(_0143_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8983_ (.D(_0144_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8984_ (.D(_0145_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8985_ (.D(_0146_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8986_ (.D(_0147_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8987_ (.D(_0148_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8988_ (.D(_0149_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8989_ (.D(_0150_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8990_ (.D(_0151_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8991_ (.D(_0152_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8992_ (.D(_0153_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8993_ (.D(_0154_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8994_ (.D(_0155_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8995_ (.D(_0156_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8996_ (.D(_0157_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8997_ (.D(_0158_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8998_ (.D(_0159_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8999_ (.D(_0160_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9000_ (.D(_0161_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9001_ (.D(_0162_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9002_ (.D(_0163_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9003_ (.D(_0164_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9004_ (.D(_0165_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9005_ (.D(_0166_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9006_ (.D(_0167_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9007_ (.D(_0168_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9008_ (.D(_0169_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9009_ (.D(_0170_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9010_ (.D(_0171_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9011_ (.D(_0172_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9012_ (.D(_0173_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9013_ (.D(_0174_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9014_ (.D(_0175_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9015_ (.D(_0176_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9016_ (.D(_0177_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9017_ (.D(_0178_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9018_ (.D(_0179_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9019_ (.D(_0180_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9020_ (.D(_0181_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9021_ (.D(_0182_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9022_ (.D(_0183_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9023_ (.D(_0184_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9024_ (.D(_0185_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9025_ (.D(_0186_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9026_ (.D(_0187_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9027_ (.D(_0188_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9028_ (.D(_0189_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9029_ (.D(_0190_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9030_ (.D(_0191_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9031_ (.D(_0192_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9032_ (.D(_0193_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9033_ (.D(_0194_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9034_ (.D(_0195_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9035_ (.D(_0196_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9036_ (.D(_0197_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9037_ (.D(_0198_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9038_ (.D(_0199_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9039_ (.D(_0200_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9040_ (.D(_0201_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9041_ (.D(_0202_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9042_ (.D(_0203_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9043_ (.D(_0204_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9044_ (.D(_0205_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9045_ (.D(_0206_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9046_ (.D(_0207_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9047_ (.D(_0208_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9048_ (.D(_0209_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9049_ (.D(_0210_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9050_ (.D(_0211_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9051_ (.D(_0212_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9052_ (.D(_0213_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9053_ (.D(_0214_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9054_ (.D(_0215_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9055_ (.D(_0216_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9056_ (.D(_0217_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9057_ (.D(_0218_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9058_ (.D(_0219_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9059_ (.D(_0220_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9060_ (.D(_0221_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9061_ (.D(_0222_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9062_ (.D(_0223_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9063_ (.D(_0224_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9064_ (.D(_0225_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9065_ (.D(_0226_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9066_ (.D(_0227_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9067_ (.D(_0228_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9068_ (.D(_0229_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9069_ (.D(_0230_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9070_ (.D(_0231_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9071_ (.D(_0232_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9072_ (.D(_0233_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9073_ (.D(_0234_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9074_ (.D(_0235_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9075_ (.D(_0236_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9076_ (.D(_0237_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9077_ (.D(_0238_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9078_ (.D(_0239_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9079_ (.D(_0240_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9080_ (.D(_0241_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9081_ (.D(_0242_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9082_ (.D(_0243_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9083_ (.D(_0244_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9084_ (.D(_0245_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9085_ (.D(_0246_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9086_ (.D(_0247_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9087_ (.D(_0248_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9088_ (.D(_0249_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9089_ (.D(_0250_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9090_ (.D(_0251_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9091_ (.D(_0252_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9092_ (.D(_0253_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9093_ (.D(_0254_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9094_ (.D(_0255_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9095_ (.D(_0256_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9096_ (.D(_0257_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9097_ (.D(_0258_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9098_ (.D(_0259_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9099_ (.D(_0260_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9100_ (.D(_0261_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9101_ (.D(_0262_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9102_ (.D(_0263_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9103_ (.D(_0264_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9104_ (.D(_0265_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9105_ (.D(_0266_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9106_ (.D(_0267_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9107_ (.D(_0268_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9108_ (.D(_0269_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9109_ (.D(_0270_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9110_ (.D(_0271_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9111_ (.D(_0272_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9112_ (.D(_0273_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9113_ (.D(_0274_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9114_ (.D(_0275_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9115_ (.D(_0276_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9116_ (.D(_0277_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9117_ (.D(_0278_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9118_ (.D(_0279_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9119_ (.D(_0280_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9120_ (.D(_0281_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9121_ (.D(_0282_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9122_ (.D(_0283_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_94 (.Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_95 (.Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9164_ (.I(net46),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9165_ (.I(net46),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9166_ (.I(net46),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9167_ (.I(net46),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9168_ (.I(net47),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9169_ (.I(net47),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9170_ (.I(net47),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(io_in[5]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(io_in[6]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[7]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input8 (.I(io_in[8]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(io_in[9]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input10 (.I(wb_rst_i),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net50),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net53),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net52),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net13),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net37),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net33),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout53 (.I(net29),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout54 (.I(net26),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_opt_3_1_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_1_wb_clk_i (.I(clknet_opt_3_0_wb_clk_i),
    .Z(clknet_opt_3_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8908__D (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8909__D (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__D (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8998__D (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9026__D (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__D (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__D (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9051__D (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9052__D (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9053__D (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__D (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__D (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__D (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9057__D (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9112__D (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9116__D (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9117__D (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9118__D (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__B (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__B2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__B (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__I (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__B (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A3 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__C (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__I (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A3 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__B1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__I (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__B2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__B2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__B (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A3 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__C (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__I (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__I (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A4 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__B (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__I (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__B2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__I (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A4 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A3 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__B (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A4 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A4 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__B1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__B1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__B (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__B (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A4 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__I0 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__B2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A3 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A3 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A3 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__I (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__I (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__B (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__B2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__B2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__I (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A4 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A4 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__I (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A4 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A4 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__C2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__B2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__I (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__B1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__B (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__B1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A3 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__C1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__C2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__B2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__B2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__B2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__B1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__I (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A4 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__B1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__B1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A2 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__B (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__I0 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__I (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__C (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__B (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__B2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__B (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__B2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__I (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__B1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__B2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__B2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__B2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A3 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__B (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__B1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__I (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A3 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__B2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__I (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__I (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__B1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__B1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__I (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__B2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__B2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__B2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__B (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A3 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A3 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A3 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A3 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__B1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__B1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__B1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__I (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__I (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__B1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__I (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__B2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__B1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A3 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__B (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__B (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__I0 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__B1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A3 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__B1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A3 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__B2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A4 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A3 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__B1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__S (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__I (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__B (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__B (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8730__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__I1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__B1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__I (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__A2 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__A2 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A2 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A2 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__C2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__B (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A2 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__B2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__B2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__B (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__I (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__B (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__I (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A2 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A3 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__B1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__B1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__B1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__C (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__I (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__I (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A3 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__B (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A3 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A4 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A4 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A3 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__B (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__C (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__C (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A3 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A3 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__B (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__C (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__C1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__C2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__B1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__B1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__B1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__B1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__I (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__B1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__C2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__I (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__C2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__B1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__B1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__I (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__I (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__I (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__C (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__C (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__C (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__B (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__C (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__C (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__B1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__B1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__C (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__A1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__C (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__C (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__B2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A4 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__C (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__C (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__B (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__C (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__B (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__B (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__C (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__B (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__I (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__C (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__B (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__B (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__B1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A2 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A2 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__B2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__B2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__B (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__C (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__B2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__B (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__B (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__B (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A2 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__B1 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__I (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__B1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__B1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__I (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__B1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__B1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__B2 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__I1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__I1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__I1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__B2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__B1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__B1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A2 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__B1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__B1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__I (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__I (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__C (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__I (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__B (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__I (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__I (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__I (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__B (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__I (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__I (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__I (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A3 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__I (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__I (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__B1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A3 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__B (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__B (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__I (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__I (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__I (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__I (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__C (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A3 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A3 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A3 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__B1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__B1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__B1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__I (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__I (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__I (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A3 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__I (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__C (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__I (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__I (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__C2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__B1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__B1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__B1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__I (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__I (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__B1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__I (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__I (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__I (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__I (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A3 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__I (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A3 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A3 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__I (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__B (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__B1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A4 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A3 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__C (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__B (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A3 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A4 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__B (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__B2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__A3 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A3 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__I (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__B2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A3 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A3 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A4 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__I (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A3 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A3 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A3 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__C (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A3 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__C (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A3 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__I (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__B2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__B2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__I (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__B2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__I (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__B2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__C (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__I (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__I (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__B (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__B (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8813__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__I (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__I (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A3 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__C (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__B (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__I (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__I (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__I (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__I (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__C (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__B (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A3 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__I (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__B (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__I (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__I (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__I (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A1 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__C (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__I (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A3 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__B (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__B2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__C (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__C (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__C (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__C (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A3 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__C (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__B (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__I (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__B (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__B (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__B (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__B (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__C2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__B (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__I (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A4 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A3 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__B2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A3 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__C (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__C (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__C (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__I (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__B (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__B (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__I (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__I (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__B2 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__B2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__B (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__C (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__B (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__I (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__I (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__B (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A3 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A2 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__I (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__B (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__C (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__B (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__B (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__B (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A3 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__I (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A4 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A3 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A3 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__I (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__C (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__C (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__B (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__B2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__I (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__I (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__I (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__I (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__I (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A1 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__I (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A3 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A4 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__I (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__I (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__I (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__I (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A3 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A4 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A3 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A3 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__I (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__B2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__I (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__I (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A4 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__B (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__I (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__B1 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A1 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A3 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A3 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__C (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A3 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__C (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__B (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__B (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__I (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A4 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__I (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__B (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A3 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__I (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A3 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A3 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A3 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__I (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__B (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__B2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__B (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A3 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A3 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__I (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__I (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__I (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__I (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__B1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__C (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A4 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__C (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A4 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__B (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__B (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__C (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__B (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__B2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__C (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__I (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__B2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A2 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__B2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__I (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__B (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__B1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__B1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__I (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__B1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__B2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__C (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__I (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__B2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8805__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__C (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__B (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__C (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A2 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A3 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A3 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__B (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__B (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__C (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__C (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__C (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__B2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__C (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A3 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A3 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A2 (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A3 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A3 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__I (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__I (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A3 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A4 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A3 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A3 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A3 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__B (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__B1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__B1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__B2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__I1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__A3 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__I (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__B (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A3 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__B (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A2 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A2 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__B (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A3 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8820__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__I1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__I1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__I (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__I (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__I (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A3 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A3 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A3 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__C (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__C (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A2 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__I (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__I (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A3 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A3 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A3 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__I (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__I (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__I (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A3 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A3 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A3 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8783__A1 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A1 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__I (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__I (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__I (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__I (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__I0 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__I (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__I (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__I (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__I (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__I (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__I (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__I (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__I (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__I (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__I (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__I (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__I (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__I (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__I (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__I (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__I0 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__I (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__I (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__I (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__I (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__I (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__I (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__I (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__C (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__C (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__I (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__I (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__I (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__I (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__B2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A1 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__I (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__I (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__I (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__I1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__C (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__C (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__I (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__I (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A3 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A3 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A3 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__I (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__I (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__B2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A2 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A3 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__C (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__C (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__C (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__I (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__S (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8821__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__I1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__S (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__S (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__S (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__S (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__B2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A3 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__I (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__I (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A4 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__B (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__I (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__I (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A4 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__I (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A3 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A3 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__I (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__C (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__I (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__B (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A3 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A3 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__I (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__C (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__I (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__C (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__I (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A2 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A2 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__B (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__B (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__B (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__C (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__C (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__I (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__B1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A2 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__I (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__A2 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A1 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A4 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__B (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A4 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__B2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__B2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A1 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__I (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A3 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__B1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__B (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__B (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A3 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__I (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A2 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A2 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A2 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__B1 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A1 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A2 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A2 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A2 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A2 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__I (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__B2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A1 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__A1 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A3 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A2 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A2 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A3 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__B2 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8717__A2 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A2 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A2 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A2 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__B1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__C (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__B1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__C (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__C (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__I (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__I (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__I (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__I (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__C (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__B (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__I (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__I (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A3 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__B (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__B (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__B (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__B (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__B (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__I (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__B (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__B (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__B (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A2 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__B (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__I0 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__C (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__C (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__I (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__I (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__I (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__B2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__B2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8755__A1 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A3 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__B1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A1 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__I (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__C (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A1 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A3 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__C (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A3 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A3 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A2 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A3 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__I (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__I (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__B2 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A3 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A3 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A4 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A3 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__I (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__I (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__B2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A3 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A3 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__I (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__C (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A4 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__B2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__I (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__I (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A4 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A1 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A3 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__B1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A1 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__C (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__B (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__I (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A2 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A3 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A3 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A3 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__I (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__I (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__S (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__S (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__S (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__S (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A2 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__I0 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__I0 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__I1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__B (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__A1 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A1 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__A1 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A1 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A1 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__B2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__I0 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A4 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A3 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A2 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__I (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__B (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__B (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A2 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__I (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A2 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A2 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A4 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A3 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__C (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A3 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A1 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__B (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__I (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__A1 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__B (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__B (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__C (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__C (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__B (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__C (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__C (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__I (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__I (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__I (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__I (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__B (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__B (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__B (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__B (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A4 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__I (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A2 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A1 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A3 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A2 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A3 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__I (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__B (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__B1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__I (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__B1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__B1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__B1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__B1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__B1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__B1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A2 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__I (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__B (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A3 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A3 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A3 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__I (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A3 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A3 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__C (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__C (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A2 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__A3 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__I (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__I (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__I (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__I (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A2 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__B (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__I (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A3 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__A3 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A2 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A2 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A3 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A2 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__B1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__C (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__A1 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__B (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__I (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A3 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A3 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__B2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__I (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__I (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__I (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__B2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__C (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A2 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__C (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__B (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__I (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__B (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A3 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__C (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__C (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__I (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__I (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A2 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__B1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__C (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A3 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__C (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A2 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__I (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__B1 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A1 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A1 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__A1 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A1 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A2 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A2 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A3 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A1 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A3 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__B (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__C (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__B (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__I (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__C (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__B (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__I (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A1 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__A1 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__B2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A1 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__I (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A2 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__C (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__C (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A2 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__B (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A4 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__B (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__I (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__I (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A1 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__C (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A2 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__B (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__I (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A1 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__B2 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__B2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__B2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__B (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__B2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__C (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__A3 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__B2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__B2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A2 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__B (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A3 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__B (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__B (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__B2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__B (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__A3 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__A2 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A1 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__B (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__I (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8826__A1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A2 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A2 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__B1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A2 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__B1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__I1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__I (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A3 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__B (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__S (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__S (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__I (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__S (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__S (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__S (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__S (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__I (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__A2 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__I1 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8837__A1 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__A1 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__I1 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__A1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__B (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8834__A1 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__B2 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__I1 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__I1 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__I1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__B (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8758__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__I (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__B (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__B (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__B (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A2 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__I (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__C (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__C (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A1 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__I (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A3 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A3 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__B1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__C (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__I (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__B (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__C (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__I (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A1 (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__C (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A2 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A2 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__B1 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__B2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__I (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__I (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__I (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__B (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A3 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__B (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__B (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A1 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__I (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A2 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A2 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A3 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A3 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A4 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__A2 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A2 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__I (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__B2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__B2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__B2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__A2 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__I (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A4 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__B (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__A2 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A1 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A2 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A2 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__C (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__I (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__B (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__B (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__C (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__B (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A3 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__C (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__B (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__B (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__B (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__A1 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A1 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A1 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__C (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A2 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A2 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__I (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__I (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A2 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A1 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A1 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__B (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__B (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A3 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__B1 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__B2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__B (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__C (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__C1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__C (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8765__I (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__C (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__C (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__B (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__B (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__C (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A2 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A2 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A3 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__B (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__B2 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__C (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A1 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A1 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A3 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__C (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A2 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__C (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__B (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__C (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__C (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__I (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__I (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__C (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__I (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__I (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__B (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__B (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A2 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__C (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__B (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__C (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A2 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__B (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8805__C (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__C (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__C (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__I (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__B2 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A2 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A2 (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__C1 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__B1 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A2 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__A2 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__A1 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__C (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__A3 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__B1 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__B2 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__C (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A3 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A1 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__A1 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__B (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__B2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__B (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__B (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A3 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A3 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__B2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__I (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A4 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__I (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__A2 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A1 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__A3 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__B (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__I (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__A2 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A2 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__I (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__A1 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__A2 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A3 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A3 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__A2 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A4 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__C (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__I (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__I (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__C (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__I (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__C (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__C (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__I (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__I (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__B2 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__B2 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__B2 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A2 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__B2 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__B2 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A2 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__I (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__B1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__B1 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A2 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A2 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__I (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__B1 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__B1 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__B1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__B1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__B1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__B1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__A2 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__B2 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A3 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A2 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A2 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__A2 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__I (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__I (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__A3 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__B (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A1 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A2 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A2 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__I (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__A2 (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__B (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A2 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A1 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A2 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__B (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__I (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__C2 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A1 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A1 (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A1 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A2 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A2 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A2 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__A2 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A2 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A2 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A2 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__B (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__B1 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__B1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__C (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A1 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__I (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__C (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__C (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__C (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__C (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__C (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A2 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A2 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A2 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A2 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A1 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A1 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__B2 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A1 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A2 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__I (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A2 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A2 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A3 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A3 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__B (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__B2 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A1 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A3 (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A2 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A1 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__B (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A2 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A2 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A2 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__B (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A2 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A3 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__B (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__C (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__C (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__C (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__B (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__A1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__I (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__A1 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A2 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A2 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__B (.I(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__C (.I(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__B (.I(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__B (.I(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A2 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7532__I (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__I (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__A2 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A1 (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__B (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A2 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__A2 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__B1 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__B2 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__C (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__C (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__B (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__C (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__A2 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A1 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__B (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__B (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__B (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A2 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A2 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A1 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A1 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__B2 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A1 (.I(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__C (.I(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__A2 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A1 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__A2 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A2 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__I (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A1 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A2 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A2 (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__B1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__I (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__B1 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__A1 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A1 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A1 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__B2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A2 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A3 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A2 (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__B1 (.I(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__B2 (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__I (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A1 (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__B2 (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__B2 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7685__A3 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A1 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A2 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A2 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A2 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__B1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__C1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__B1 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A2 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A2 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__B2 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__B2 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A1 (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A1 (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A1 (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A2 (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__A2 (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__B1 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A1 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A1 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A2 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A3 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__A2 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A2 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A1 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A2 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A2 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__I (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A2 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A2 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A2 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__I (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A1 (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__A1 (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A2 (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A1 (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A3 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__B (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__B1 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A1 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A1 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__C (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__B (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__B (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__B2 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A2 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A2 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__A1 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__B2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__B2 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A1 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A1 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__B (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__C (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A2 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__I (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A1 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A1 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__B (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__C1 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__B1 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__I (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__A1 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A1 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__B2 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__B2 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__B (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A1 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__B (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__B (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__I (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__B (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__I (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A1 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A1 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A1 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__I (.I(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A2 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A2 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A2 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A3 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A2 (.I(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__A1 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__B2 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__B (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__B (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__B (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__B (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__B2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__B (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__B (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A2 (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A1 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A1 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__B (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A1 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__A1 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A1 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A1 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__B (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A2 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8454__A1 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A3 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__B (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__B1 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__B1 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__B1 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__B1 (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__B1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A2 (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__B1 (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__B2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__A2 (.I(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A1 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__B1 (.I(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A2 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A1 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__B (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A2 (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__A2 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A2 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A2 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A2 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A2 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__B (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A3 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__B2 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__B (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A1 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__B1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__B (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A2 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A1 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A3 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__B1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A3 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__B2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__B2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A2 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A1 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A1 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A3 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__B (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__B1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A1 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__I (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__C (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A1 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A1 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__B2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A1 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A1 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A1 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__C (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__A2 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__C (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__B (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__B (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__B (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__B (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__B (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A1 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__A1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__I (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__A1 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A1 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__B1 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__B2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__B2 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__B1 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A2 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__A1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__A1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__B (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A2 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__B (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__C (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__B2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__B1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__I (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A2 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__B1 (.I(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A2 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A2 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A2 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__B (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__C (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A2 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A4 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__I (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__A3 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A2 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__A2 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__A2 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A2 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A2 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A2 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__A1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__B (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A2 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__A2 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__B (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__B1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__B2 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A4 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A3 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A2 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A2 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__B1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__B1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__A2 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__B1 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__A4 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A2 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__C (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__B (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__A2 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__B1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__B (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A2 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A2 (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__B (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__B (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__B (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__B (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__B (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__B1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__B1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__A2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__B (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__C (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__A2 (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__B1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__B (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__B2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__B1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__B (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A2 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__A1 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A1 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A3 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A3 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A4 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A3 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__B (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__B (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__B (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__C (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__C (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__S (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__S (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__I (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__B (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__I (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__I (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A3 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__I (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A2 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__B1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__B1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__B1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__C (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__B (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__A2 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A2 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__B1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A2 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__C1 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__B1 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A3 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__C (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__B (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__I (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__I (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__B (.I(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__B (.I(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__B (.I(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__B (.I(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A1 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A1 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__C (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__C (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__B2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__B (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__B (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A2 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A2 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__B1 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__B (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__B2 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__I (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8758__A2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__C (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__C (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A1 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__C (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__B2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__C (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__B (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__C (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__A1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__B (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__B1 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__B (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__B2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__B (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__B1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__C (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A1 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__B (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A1 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__B (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__B1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__C (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__B (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__B (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__A1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__B1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__B (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A1 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A1 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A1 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A1 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A2 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__A1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__A1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__B (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__B1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__B2 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__B (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__I0 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__B (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__B1 (.I(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__C (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__I0 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__A1 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__B (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A3 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__B (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__I (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__I (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__B1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__B1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__B1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__C (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__C (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__I (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__I (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__C (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__C (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__I (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__I (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__I (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A2 (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A2 (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A2 (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__I (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__A2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__A2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__I (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__I (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A2 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A2 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__I (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__I (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A2 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A2 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A2 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A2 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A3 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__B (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__B2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__B2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__A1 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A1 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A1 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__B (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__B (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__A1 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A1 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A2 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A1 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__B (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A1 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__I (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A1 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__B1 (.I(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__B1 (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__B (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A1 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__B2 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__C (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__I (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__C (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__B2 (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__I (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__I (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__I (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A2 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A2 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__A2 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__B1 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A2 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__I (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__I (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A2 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A2 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A2 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__B1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__B (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__C (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__C (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__C (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__B1 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__B (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__B1 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__B1 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A2 (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A2 (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__B2 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A2 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__A1 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__I (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__B (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A2 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A2 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A1 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__B (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__B (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__B (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__B (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A2 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A2 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A2 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A2 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__B1 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A2 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__B1 (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A2 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__B (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__B2 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__B1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__B1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A2 (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__C (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__A2 (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A2 (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A2 (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__A2 (.I(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__B (.I(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A2 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A2 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A3 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A2 (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__B (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A2 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__A1 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__B (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__B (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__B (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__B (.I(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A1 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__A2 (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__B2 (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__B (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__A1 (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__A1 (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__A1 (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A1 (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__A2 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A2 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__B1 (.I(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__B2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__A1 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A1 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__B2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A1 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A1 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A2 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A1 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A2 (.I(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__C (.I(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__B (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__B1 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__B (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A1 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__C (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__C (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A1 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A2 (.I(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A2 (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A2 (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__B (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A3 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A2 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__B (.I(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__B (.I(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__B1 (.I(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__B2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__B2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__B2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__B2 (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__C (.I(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8823__C (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__C (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__C (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__C (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__B2 (.I(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A1 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__A1 (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A1 (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A1 (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A1 (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__B (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A2 (.I(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__B1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__C (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__B (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A1 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A2 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A1 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__B1 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__C (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__B (.I(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__A1 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A2 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A1 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A2 (.I(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A2 (.I(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__A1 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__A2 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__A1 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A2 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__B1 (.I(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A2 (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__A2 (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__A2 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__A2 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__A2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__B1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__B (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__B1 (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__B2 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A1 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A3 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A4 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A3 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A2 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__A2 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A1 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__B2 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A1 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A2 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__B1 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A2 (.I(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__B1 (.I(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__A2 (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A2 (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__B1 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__I (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__I (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__A2 (.I(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__A2 (.I(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__A2 (.I(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__A2 (.I(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__A2 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__A2 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__A2 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__A2 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__A2 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A2 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__A2 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__A2 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__A3 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__I (.I(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__A2 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__A1 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A1 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__A2 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A2 (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__A2 (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__B (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__B (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__B (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__A2 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__A2 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__A2 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__A2 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__B (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__A2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__A1 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__A1 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__A1 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__A1 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__A2 (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__B (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__A2 (.I(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__B (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__A2 (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A1 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__C (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__A1 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__A1 (.I(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__A3 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__A1 (.I(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__A1 (.I(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__B (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__A2 (.I(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__B (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__A1 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__A2 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__A2 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__A2 (.I(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__A1 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8820__A3 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8801__A1 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__A1 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__A2 (.I(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A2 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__B (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__B2 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__A2 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A2 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A2 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__A2 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8762__A1 (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__A2 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__A1 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A1 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A3 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A2 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__A2 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8783__A2 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__A1 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__A2 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__A1 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A1 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__A2 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A2 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__A2 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8805__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__B (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8805__B2 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__B (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A2 (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__A3 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8813__A2 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A3 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8823__A1 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8822__A2 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__B (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__B (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__C (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8826__B (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8827__I (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__I (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__C (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__S0 (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__S0 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__S0 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__I (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__A1 (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A1 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A1 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__I (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__I (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__I (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__S (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__S (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__S (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__I (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S1 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__S (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__S (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__S (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__S1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__S (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__S (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__I (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__S1 (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__B2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__S0 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__S0 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__S0 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__I (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__I (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__S1 (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A2 (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A1 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A1 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__I (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A2 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__I (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__I (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A4 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__I (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__I (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__I (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__I (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__I (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__I (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__I (.I(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A1 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__I (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A3 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A1 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__I (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A2 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__A1 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__A4 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__I (.I(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A1 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A2 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A2 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A3 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__B (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__I (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A2 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A4 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A1 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__I (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A3 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A3 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A2 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__I (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A3 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__I (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__B (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__I (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A1 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A2 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A2 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__I (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__I (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A2 (.I(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A2 (.I(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__I (.I(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A3 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A1 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__I (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__I (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A1 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A1 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__B (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__I (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__I (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A1 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A1 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A1 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A1 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A2 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__B2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A2 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__A1 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__I (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__B (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A3 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A2 (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__B (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__I (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A2 (.I(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A3 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A2 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A3 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__I (.I(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A1 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__I (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__I (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A3 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A2 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A3 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A2 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__I (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A1 (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A2 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__I (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A2 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__I (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__I (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A2 (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A2 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A3 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__I (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A3 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A3 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A1 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A2 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__A2 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__A2 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A4 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A2 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__I (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A1 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A3 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__I (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__C (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__I (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A3 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A1 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__I (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__I (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__I (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A3 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__B (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__S (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__C (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I0 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__I (.I(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I1 (.I(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I3 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__B (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__I (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__I1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__I (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__S (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A2 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__I (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A2 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A2 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__B (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A1 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__B (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__B (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__C (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__B (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A1 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__I (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A2 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__I (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__B2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__B1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__B (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__I (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__B (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__A1 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__B (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__B (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__A2 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A1 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A3 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__I (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__B2 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__I (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__I (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__I (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A2 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A1 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A1 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A1 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__I (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__B3 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__C (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__C (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__I (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__I (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A3 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__C (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__I (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__I (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__C (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__C (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__C (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__I (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__B2 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__I (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__A1 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__B2 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A1 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A1 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A1 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__I (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__B2 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__I (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__I (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A3 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A1 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__I (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__B1 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__I (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__I (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__C (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__I (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__I (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__B2 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__I (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A1 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__I (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A1 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A3 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A4 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A3 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A3 (.I(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__S (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A2 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A1 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A1 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__I (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A1 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__C2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__I (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A1 (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__I (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__I (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__I (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__I (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A2 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__I (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__B (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A1 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__C (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__B (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__B (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__C (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__B (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__A1 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A1 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A1 (.I(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__B (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A2 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__I (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A2 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A2 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A2 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__B (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__I (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__B (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__I (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__B (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A2 (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A2 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A2 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__B1 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A1 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__C (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__I (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__I (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__C (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A1 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A1 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__I (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__I (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__I (.I(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A2 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__B (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__I (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A1 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A2 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__B (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__I (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__I (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__I (.I(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A1 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__I (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A2 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A2 (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__I (.I(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__C (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__I (.I(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__B2 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__I (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A3 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A3 (.I(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A1 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A1 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A2 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A3 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A1 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A1 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I1 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A1 (.I(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A1 (.I(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I (.I(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__I (.I(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__A1 (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__A2 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A3 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A1 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A2 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__I (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__I (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__B2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__B2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__B2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__I (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__I (.I(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A3 (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__I (.I(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A2 (.I(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A3 (.I(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A1 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A2 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A2 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A3 (.I(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A1 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A1 (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__I (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A3 (.I(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A1 (.I(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A2 (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A4 (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__B2 (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__B (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__B1 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__C (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__C (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A3 (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A4 (.I(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__A2 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A2 (.I(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A1 (.I(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A2 (.I(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__B (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__B2 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A2 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A2 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A1 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__I (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A1 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A1 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A1 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__A1 (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__I (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A3 (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A1 (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__C (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__I (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__I (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__B (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__B2 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A2 (.I(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A2 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A2 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__B2 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A2 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__I (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__I (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A1 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__I (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A2 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A1 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A1 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A3 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__I (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__B1 (.I(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__I (.I(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__I (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A3 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A2 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A1 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A1 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A1 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__I (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A1 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__I (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__I (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__C1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A2 (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__B (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A2 (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A2 (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A3 (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A2 (.I(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__B (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A3 (.I(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A2 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A2 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A2 (.I(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A2 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A2 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__I (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__I (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A4 (.I(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__B1 (.I(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__I (.I(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A1 (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A2 (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__B1 (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A4 (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A1 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__B2 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A1 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__I (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A1 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A1 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A1 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__I (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__I (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__I0 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__I0 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A1 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__I (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__I (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__I (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A3 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A2 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A2 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A1 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A1 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8822__B (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__I (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__I (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__I (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8836__B (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__I (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__I (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I0 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__I (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__I (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I0 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I0 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I0 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I0 (.I(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I0 (.I(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I0 (.I(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B2 (.I(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I0 (.I(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__B2 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__B2 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__I1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I3 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__B2 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__I1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I3 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__A1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__B2 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__B2 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__B2 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__I1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__B2 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I3 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I1 (.I(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A1 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I2 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__B2 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__A1 (.I(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__B2 (.I(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__B2 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__B2 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__B2 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__B2 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__C1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__I1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__B2 (.I(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__B2 (.I(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__B2 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__B2 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__I1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__B2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__B2 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__B2 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__B2 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__B2 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__B2 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__B2 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__B2 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__B2 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__B2 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__B2 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__B2 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__B2 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__C1 (.I(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__B2 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__B2 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__B2 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__B2 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__B2 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__B2 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__B2 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__B2 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__B2 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__B2 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A1 (.I(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A1 (.I(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A1 (.I(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__B2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A3 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9167__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9166__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9165__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9164__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__B2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8968__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8985__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9018__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9017__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9021__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9022__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9109__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8910__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8913__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8912__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9110__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9106__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9105__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9104__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9102__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9103__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9101__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9014__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9002__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9028__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9029__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9027__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9026__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9032__CLK (.I(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9090__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9085__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9083__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9081__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9084__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9082__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9091__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9093__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9086__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9088__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9089__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9087__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9092__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9045__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9044__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9043__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8924__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9037__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8923__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8920__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8926__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8928__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8929__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8946__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8917__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8914__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8916__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8919__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8947__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8950__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8949__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8948__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8915__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8972__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8973__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9063__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8941__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8939__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8943__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9061__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9062__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9069__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9073__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9067__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9058__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9048__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9060__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9064__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8927__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9036__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9046__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9065__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9059__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9072__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8890__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9070__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9111__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8938__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8940__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9115__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9066__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9071__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9068__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9113__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8960__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8955__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8942__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9119__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9116__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9121__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8882__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8868__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8875__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8874__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8861__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9118__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8855__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8959__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8954__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8880__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8958__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9112__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8860__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8881__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9098__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8873__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8859__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8867__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8869__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8887__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9078__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9074__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9094__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8883__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8896__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8885__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9077__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8894__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8884__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8892__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9076__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9096__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8864__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8863__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9075__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9097__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8871__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8856__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9095__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8961__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8956__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8944__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8870__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8857__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8976__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8977__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8858__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8865__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8951__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8952__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8953__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8975__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8905__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8906__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8889__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8851__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9057__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9117__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9052__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9051__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8849__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8989__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8850__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8991__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8990__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8854__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8852__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8993__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8844__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8846__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8988__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8986__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8965__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8964__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9007__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9008__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8978__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8963__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8962__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8848__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9023__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9003__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9025__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8998__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9031__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8899__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8931__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8898__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9120__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9039__CLK (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8901__CLK (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__CLK (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_1_wb_clk_i_I (.I(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_opt_3_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net90;
 assign io_oeb[13] = net95;
 assign io_oeb[14] = net55;
 assign io_oeb[15] = net56;
 assign io_oeb[16] = net57;
 assign io_oeb[17] = net58;
 assign io_oeb[18] = net59;
 assign io_oeb[19] = net60;
 assign io_oeb[1] = net91;
 assign io_oeb[20] = net61;
 assign io_oeb[21] = net62;
 assign io_oeb[22] = net63;
 assign io_oeb[23] = net64;
 assign io_oeb[24] = net65;
 assign io_oeb[25] = net66;
 assign io_oeb[26] = net67;
 assign io_oeb[27] = net68;
 assign io_oeb[28] = net69;
 assign io_oeb[29] = net70;
 assign io_oeb[2] = net92;
 assign io_oeb[30] = net71;
 assign io_oeb[31] = net72;
 assign io_oeb[32] = net73;
 assign io_oeb[33] = net74;
 assign io_oeb[34] = net75;
 assign io_oeb[35] = net76;
 assign io_oeb[36] = net77;
 assign io_oeb[37] = net78;
 assign io_oeb[3] = net93;
 assign io_oeb[4] = net94;
 assign io_out[0] = net79;
 assign io_out[13] = net84;
 assign io_out[1] = net80;
 assign io_out[2] = net81;
 assign io_out[33] = net85;
 assign io_out[34] = net86;
 assign io_out[35] = net87;
 assign io_out[36] = net88;
 assign io_out[37] = net89;
 assign io_out[3] = net82;
 assign io_out[4] = net83;
endmodule

