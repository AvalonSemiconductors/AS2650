* NGSPICE file created from gpios.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

.subckt gpios DAC_clk DAC_d1 DAC_d2 DAC_le RXD TXD addr[0] addr[1] addr[2] addr[3]
+ bus_cyc bus_we data_in[0] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5]
+ data_in[6] data_in[7] data_out[0] data_out[1] data_out[2] data_out[3] data_out[4]
+ data_out[5] data_out[6] data_out[7] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] irq0 irq6 irq7 la_data_out[0] la_data_out[1] la_data_out[2]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] pwm0
+ pwm1 pwm2 rst tmr0_clk tmr0_o tmr1_clk tmr1_o vdd vss wb_clk_i
XTAP_TAPCELL_ROW_52_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_432_ PORTB\[2\] _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_501_ _134_ _114_ _125_ _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_23_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__568__A1 DDRB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__568__B2 DDRA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__740__A1 PORTA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_415_ _078_ net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__789__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__713__A1 _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input36_I pwm0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__704__A1 DDRB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_895_ _060_ clknet_3_6__leaf_wb_clk_i SPB\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_680_ _258_ _279_ _288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_878_ _043_ clknet_3_7__leaf_wb_clk_i PORTA\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__844__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_732_ _248_ _326_ _327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__867__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_801_ SPA\[6\] _370_ _378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_7__f_wb_clk_i clknet_0_wb_clk_i clknet_3_7__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_594_ _218_ _120_ _213_ _219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_663_ net15 _275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__437__I0 PORTB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__786__B _359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput75 net75 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 net42 RXD vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput64 net64 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput53 net53 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_715_ _227_ _313_ _314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput86 net99 la_data_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_577_ _202_ _203_ _149_ _101_ _204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__595__A2 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_646_ _261_ _262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__535__I _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_500_ _107_ _134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_48_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_431_ SPB\[2\] _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_8_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_629_ net16 _248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_46_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__495__A1 DDRB\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_414_ PORTA\[6\] net37 SPA\[6\] _078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_19_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__713__A2 _263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input29_I io_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__401__A1 _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_894_ _059_ clknet_3_6__leaf_wb_clk_i SPA\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__622__A1 _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_6__f_wb_clk_i clknet_0_wb_clk_i clknet_3_6__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_877_ _042_ clknet_3_7__leaf_wb_clk_i PORTA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_731_ _312_ _326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_662_ _273_ _274_ _262_ _022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_800_ _218_ _364_ _377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_593_ net18 _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__834__A1 _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__696__C _254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__825__A1 SPB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput76 net76 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput87 net97 la_data_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput65 net65 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput54 net54 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput43 net43 data_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_714_ _312_ _313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_645_ net39 _261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_576_ _113_ _121_ _130_ _141_ _203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_41_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I DAC_d2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__807__A1 _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__857__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_430_ _084_ net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__461__I _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_628_ _246_ _236_ _247_ _241_ _015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_559_ net48 _188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__495__A2 _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_413_ _077_ net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_5__f_wb_clk_i clknet_0_wb_clk_i clknet_3_5__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_893_ _058_ clknet_3_2__leaf_wb_clk_i SPA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_43_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input41_I tmr1_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_876_ _041_ clknet_3_7__leaf_wb_clk_i PORTA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__890__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_730_ _324_ _325_ _323_ _039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_592_ _099_ _217_ _009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_661_ DDRA\[2\] _268_ _274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__464__I _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_859_ _024_ clknet_3_0__leaf_wb_clk_i DDRA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__770__A1 _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput77 net77 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput88 net100 la_data_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput66 net66 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput55 net55 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 net44 data_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_575_ net26 _202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_644_ net93 _244_ _260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_713_ _135_ _263_ _312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__743__A1 _258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__734__A1 PORTA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_627_ net15 _235_ _247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_558_ _171_ _180_ _184_ _187_ _170_ _005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_13_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_489_ _122_ _123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_14_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_4__f_wb_clk_i clknet_0_wb_clk_i clknet_3_4__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_412_ PORTA\[5\] net36 SPA\[5\] _077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__707__A1 DDRB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__472__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__847__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_892_ _057_ clknet_3_2__leaf_wb_clk_i SPA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__467__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input34_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_875_ _040_ clknet_3_7__leaf_wb_clk_i PORTA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__534__C1 SPA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_591_ net83 _214_ _216_ _217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_660_ _242_ _265_ _273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_51_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__480__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_858_ _023_ clknet_3_0__leaf_wb_clk_i DDRA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_789_ net15 _365_ _369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__589__A2 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput78 net78 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput67 net67 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput89 net98 la_data_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output65_I net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput56 net56 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_712_ _310_ _311_ _309_ _035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput45 net45 data_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_643_ _258_ _230_ _259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_574_ net50 _201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__880__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_3__f_wb_clk_i clknet_0_wb_clk_i clknet_3_3__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_626_ net89 _246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_557_ _185_ _186_ _187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__422__A1 SPA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_488_ _113_ _121_ _117_ _118_ _122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_14_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__661__A1 DDRA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__716__A2 _263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_411_ _076_ net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__643__A1 _258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_609_ _227_ _231_ _232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__663__I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__634__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_891_ _056_ clknet_3_2__leaf_wb_clk_i SPA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_16_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input27_I io_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__837__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_874_ _039_ clknet_3_7__leaf_wb_clk_i PORTA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__478__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__828__A1 SPB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_590_ last_irq0_trigger _215_ _216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__819__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_788_ _073_ _362_ _368_ _346_ _054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_3_2__f_wb_clk_i clknet_0_wb_clk_i clknet_3_2__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_857_ _022_ clknet_3_1__leaf_wb_clk_i DDRA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput57 net57 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__514__C _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput46 net46 data_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput68 net68 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput79 net79 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_711_ DDRB\[7\] _302_ _311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_642_ net19 _258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_573_ _171_ _195_ _196_ _200_ _098_ _007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_625_ _243_ _245_ _238_ _014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__422__A2 DDRA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_556_ SPB\[4\] _111_ _163_ net23 _144_ _186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_487_ _108_ _121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I DAC_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__870__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__652__A2 _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_410_ PORTA\[4\] net41 SPA\[4\] _076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__702__C _254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_608_ _230_ _231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_19_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_539_ _104_ _158_ _162_ _169_ _170_ _003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_27_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__893__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__570__A1 SPB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_890_ _055_ clknet_3_2__leaf_wb_clk_i SPA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_16_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__561__A1 _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__584__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__791__A1 SPA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_873_ _038_ clknet_3_5__leaf_wb_clk_i PORTA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_3_1__f_wb_clk_i clknet_0_wb_clk_i clknet_3_1__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__494__I _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__782__A1 _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__534__A1 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__773__A1 _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_787_ net14 _361_ _368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_856_ _021_ clknet_3_1__leaf_wb_clk_i DDRA\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__620__C _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__746__A1 _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput69 net69 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_43_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput47 net47 data_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput58 net58 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_641_ _256_ _257_ _238_ _018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_572_ _197_ _198_ _199_ _200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_710_ _258_ _291_ _310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__737__A1 PORTA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_839_ _004_ clknet_3_4__leaf_wb_clk_i net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__728__A1 _275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__525__C _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_624_ net88 _244_ _245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_48_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_555_ net90 _133_ _167_ PORTA\[4\] SPA\[4\] _165_ _185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_54_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_486_ _119_ _120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__412__I0 PORTA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__497__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_538_ _097_ _170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_607_ _228_ _229_ _230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_469_ _102_ _103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__555__C1 SPA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0__f_wb_clk_i clknet_0_wb_clk_i clknet_3_0__leaf_wb_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_16_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__860__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_872_ _037_ clknet_3_5__leaf_wb_clk_i PORTA\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__883__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__519__C1 SPA\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__782__A2 _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input32_I io_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__719__B _309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_855_ _020_ clknet_3_1__leaf_wb_clk_i DDRA\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_786_ _366_ _367_ _359_ _053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_27_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__746__A2 _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput48 net48 data_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput59 net59 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_640_ net92 _244_ _257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_571_ PORTB\[6\] _128_ _119_ net84 _199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__425__A1 SPA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_838_ _003_ clknet_3_1__leaf_wb_clk_i net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_769_ _353_ _354_ _349_ _049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__664__A1 _275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_623_ _234_ _244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_554_ PORTB\[4\] _155_ _174_ DDRA\[4\] _183_ _184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_485_ _113_ _115_ _117_ _118_ _119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_54_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__412__I1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__403__I1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_468_ _101_ _102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_537_ _166_ _168_ _169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__800__A1 _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_606_ _101_ net11 _229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__555__B1 _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__412__S SPA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_871_ _036_ clknet_3_5__leaf_wb_clk_i PORTA\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input25_I io_in[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_854_ _019_ clknet_3_5__leaf_wb_clk_i net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__850__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_785_ SPA\[1\] _362_ _367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__873__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput49 net49 data_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_54_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_570_ SPB\[6\] _154_ _163_ net25 _144_ _198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__425__A2 _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_768_ PORTB\[5\] _351_ _354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_837_ _002_ clknet_3_1__leaf_wb_clk_i net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_699_ DDRB\[3\] _302_ _303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__896__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_622_ _242_ _231_ _243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_484_ net9 _118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_553_ _181_ _159_ _160_ _182_ _183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__591__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_605_ _134_ _115_ _117_ _118_ _228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_54_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__564__A1 SPB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__564__B2 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_536_ PORTA\[2\] _167_ _143_ DDRA\[2\] _103_ _168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_467_ net10 _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__637__C _254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__555__B2 PORTA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__546__A1 PORTB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__794__A1 SPA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__785__A1 SPA\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_519_ net35 _140_ _136_ PORTA\[1\] SPA\[1\] _138_ _152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_15_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_21_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_870_ _035_ clknet_3_1__leaf_wb_clk_i DDRB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__767__A1 _283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__758__A1 _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input18_I data_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__749__A1 _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_853_ _018_ clknet_3_4__leaf_wb_clk_i net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_784_ _270_ _365_ _366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_767_ _283_ _337_ _353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_836_ _001_ clknet_3_1__leaf_wb_clk_i net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_698_ _294_ _302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__840__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_621_ net14 _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_54_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_552_ net30 _182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_483_ _116_ _117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__863__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_819_ net16 _384_ _390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__405__I SPA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__886__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_535_ _135_ _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_604_ net12 _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_466_ _099_ _100_ _000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__491__A1 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__901__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_518_ _149_ _150_ _151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_51_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_449_ SPB\[7\] DDRB\[7\] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__519__A2 _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__455__A1 _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__446__A1 SPB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__659__B _262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_852_ _017_ clknet_3_5__leaf_wb_clk_i net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_783_ _364_ _365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__600__A1 _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input30_I io_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__419__A1 SPA\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_904_ _069_ clknet_3_6__leaf_wb_clk_i last_irg6_trigger vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_766_ _350_ _352_ _349_ _048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_835_ _000_ clknet_3_6__leaf_wb_clk_i last_irq7_trigger vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_697_ _275_ _292_ _301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__830__A1 _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__821__A1 SPB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__429__S SPB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_620_ _239_ _236_ _240_ _241_ _013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_551_ DDRB\[4\] _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__812__A1 SPB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_482_ net8 _116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_818_ _087_ _381_ _389_ _147_ _063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_54_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__803__A1 _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_749_ _127_ _212_ _340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_534_ net21 _163_ _164_ net88 SPA\[2\] _165_ _166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_465_ SPA\[7\] net33 _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_603_ _099_ _226_ _011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_54_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__416__I SPA\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__853__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_448_ SPB\[6\] DDRB\[6\] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_517_ DDRB\[1\] _126_ _143_ DDRA\[1\] _150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__437__S SPB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__876__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__455__A2 _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__899__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_851_ _016_ clknet_3_5__leaf_wb_clk_i net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_782_ _137_ _233_ _364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_32_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__604__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input23_I io_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_903_ _068_ clknet_3_7__leaf_wb_clk_i last_irq0_trigger vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_834_ _241_ _220_ _069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_765_ PORTB\[4\] _351_ _352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__594__A1 _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_696_ _093_ _296_ _300_ _254_ _030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_6_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__649__A2 _263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__585__A1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_550_ net47 _180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_481_ _114_ _115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_32_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_817_ net15 _380_ _389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_748_ _210_ _338_ _339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_679_ _286_ _287_ _278_ _026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__577__C _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_602_ net85 _224_ _225_ _226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__797__A1 SPA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_533_ _137_ _165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_464_ _098_ _099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__788__A1 _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__522__I _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__703__A1 _283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_35_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_447_ SPB\[5\] DDRB\[5\] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_15_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_516_ _121_ _130_ _118_ _149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_50_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__843__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_850_ _015_ clknet_3_5__leaf_wb_clk_i net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_781_ _070_ _362_ _363_ _346_ _052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__776__B _359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__866__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__600__A3 _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input16_I data_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output84_I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_833_ _241_ _215_ _068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__889__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_764_ _340_ _351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_902_ _067_ clknet_3_3__leaf_wb_clk_i SPB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_695_ net14 _295_ _300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__615__I _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input8_I addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__585__A2 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_480_ net7 _114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_22_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_747_ _337_ _338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_816_ _387_ _388_ _376_ _062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__904__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_678_ DDRA\[6\] _281_ _287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_601_ last_irq7_trigger _100_ _225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_4_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_532_ _132_ _164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_463_ _097_ _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_515_ net44 _148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_446_ SPB\[4\] DDRB\[4\] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__458__A1 _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__630__A1 _248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__533__I _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__697__A1 _275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__449__A1 SPB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_429_ PORTB\[1\] net38 SPB\[1\] _084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 DAC_clk net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_780_ _210_ _361_ _363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__833__A1 _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__792__B _359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__824__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_901_ _066_ clknet_3_3__leaf_wb_clk_i SPB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_763_ _248_ _338_ _350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_694_ _298_ _296_ _299_ _254_ _029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__815__A1 _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_832_ _398_ _399_ _393_ _067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__594__A3 _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__856__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_746_ _127_ _233_ _337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_677_ _255_ _279_ _286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_815_ _085_ _381_ _388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__879__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_531_ _140_ _163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_600_ _223_ _120_ _213_ _224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_4_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_462_ net39 _097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_729_ PORTA\[3\] _316_ _325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__694__C _254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_514_ _104_ _105_ _124_ _146_ _147_ _001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_51_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_445_ SPB\[1\] DDRB\[1\] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__458__A2 net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__795__B _359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input39_I rst vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__449__A2 DDRB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_428_ _083_ net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput2 DAC_d1 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__597__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__629__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__588__A1 _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__760__A1 PORTB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_900_ _065_ clknet_3_3__leaf_wb_clk_i SPB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_831_ SPB\[7\] _391_ _399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__579__B2 SPA\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_762_ _347_ _348_ _349_ _047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_693_ net13 _295_ _299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input21_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_814_ _242_ _384_ _387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_745_ _335_ _336_ _334_ _043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_676_ _284_ _285_ _278_ _025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__724__A1 PORTA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__642__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__715__A1 _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_461_ _096_ net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_530_ SPB\[2\] _111_ _155_ PORTB\[2\] _161_ _162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_54_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__462__I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__706__A1 _255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_728_ _275_ _313_ _324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_659_ _271_ _272_ _262_ _021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_1_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__846__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_444_ _092_ net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_513_ _097_ _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__869__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_427_ _082_ PORTB\[0\] _083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_15_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__439__I0 PORTB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 DAC_d2 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__645__I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_761_ _322_ _349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_830_ _223_ _383_ _398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_692_ DDRB\[1\] _298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_26_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_10_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input14_I data_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_744_ PORTA\[7\] _328_ _336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_813_ _385_ _386_ _376_ _061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__421__A1 SPA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_675_ DDRA\[5\] _281_ _285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input6_I addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__660__A1 _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__651__A1 _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_460_ SPB\[3\] net22 _096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_727_ _320_ _321_ _323_ _038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_589_ SPA\[0\] net20 _215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_658_ DDRA\[1\] _268_ _272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_443_ PORTB\[7\] net1 SPB\[7\] _092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_512_ _129_ _139_ _145_ _146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__473__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__560__C2 PORTB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__606__A1 _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__468__I _101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_426_ SPB\[0\] _082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_11_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__836__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 DAC_le net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_40_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__827__A1 _218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__859__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_409_ _075_ net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__809__A1 _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__588__A3 _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_760_ PORTB\[3\] _341_ _348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_691_ _293_ _297_ _290_ _028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__656__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_889_ _054_ clknet_3_7__leaf_wb_clk_i SPA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput40 tmr0_o net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_743_ _258_ _326_ _335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_674_ _283_ _279_ _284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_812_ SPB\[1\] _381_ _386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__421__A2 DDRA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_726_ _322_ _323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_657_ _270_ _265_ _271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_588_ _210_ _120_ _213_ _214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_39_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__892__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_511_ net34 _140_ _143_ DDRA\[0\] _144_ _145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_442_ _091_ net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__560__B2 DDRA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__560__A1 DDRB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_709_ _307_ _308_ _309_ _034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__606__A2 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__484__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_425_ SPA\[2\] _081_ net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__781__A1 _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 TXD net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input37_I pwm1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__763__A1 _248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_408_ PORTA\[3\] net40 SPA\[3\] _075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__809__A2 _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_690_ DDRB\[0\] _296_ _297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__736__A1 _283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_888_ _053_ clknet_3_3__leaf_wb_clk_i SPA\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_16_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput30 io_in[4] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 tmr1_o net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__849__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_811_ net13 _384_ _385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_742_ _332_ _333_ _334_ _042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_673_ net17 _283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_53_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__581__C1 _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_656_ net13 _270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_725_ net39 _322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_587_ _212_ _213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_441_ PORTB\[6\] net4 SPB\[6\] _091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_510_ _102_ _144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__545__C1 SPA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_639_ _255_ _231_ _256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_708_ _261_ _309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_424_ net28 _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__882__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 addr[0] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__460__A1 SPB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__451__A1 _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__709__B _309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_407_ _074_ net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__690__A1 DDRB\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__433__A1 _085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_887_ _052_ clknet_3_7__leaf_wb_clk_i SPA\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput31 io_in[5] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 io_in[0] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__654__A1 DDRA\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_810_ _383_ _384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__406__A1 _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_741_ _322_ _334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_672_ _280_ _282_ _278_ _024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__722__B _309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input12_I data_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__593__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_724_ PORTA\[2\] _316_ _321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__627__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_655_ _266_ _269_ _262_ _020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_18_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_586_ _211_ _212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_26_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__839__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__618__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I DAC_le vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__609__A1 _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_440_ _090_ net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__545__B1 _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_707_ DDRB\[6\] _302_ _308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_569_ net92 _133_ _136_ PORTA\[6\] SPA\[6\] _138_ _197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_638_ net18 _255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_37_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_423_ SPA\[6\] DDRA\[6\] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 addr[1] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__451__A2 DDRA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_406_ _073_ PORTA\[2\] _074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_28_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_44_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__433__A2 _086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__872__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_886_ _051_ clknet_3_6__leaf_wb_clk_i PORTB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput21 io_in[10] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput32 io_in[6] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 bus_cyc net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__410__S SPA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__895__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_740_ PORTA\[6\] _328_ _333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_7_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__406__A2 PORTA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_671_ DDRA\[4\] _281_ _282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_5_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_869_ _034_ clknet_3_2__leaf_wb_clk_i DDRB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__581__A1 SPB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__581__B2 PORTB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_723_ _242_ _313_ _320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_31_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_654_ DDRA\[0\] _268_ _269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_585_ net10 net11 _211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_26_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__563__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__554__B2 DDRA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__554__A1 PORTB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__490__C2 net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__793__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__545__B2 PORTA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_637_ _251_ _236_ _252_ _254_ _017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_706_ _255_ _292_ _307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_499_ _132_ _133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__536__B2 DDRA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__536__A1 PORTA\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_568_ DDRB\[6\] _173_ _174_ DDRA\[6\] _123_ net32 _196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__784__A1 _270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__599__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_422_ SPA\[5\] DDRA\[5\] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_11_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 addr[2] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_52_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__748__A1 _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__739__A1 _255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_405_ SPA\[2\] _073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_51_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__408__S SPA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input35_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__441__I0 PORTB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_885_ _050_ clknet_3_6__leaf_wb_clk_i PORTB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput22 io_in[11] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 io_in[7] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput11 bus_we net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_670_ _267_ _281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__414__I0 PORTA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_868_ _033_ clknet_3_2__leaf_wb_clk_i DDRB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_799_ _374_ _375_ _376_ _057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__862__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_722_ _318_ _319_ _309_ _037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_653_ _267_ _268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_18_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_584_ net12 _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__885__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__490__B2 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__818__C _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__545__A2 _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_567_ net49 _195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_705_ _305_ _306_ _290_ _033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_636_ _253_ _254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__536__A2 _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_498_ _112_ _108_ _130_ _131_ _132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_41_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__900__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_421_ SPA\[4\] DDRA\[4\] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_11_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 addr[3] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_619_ _097_ _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__693__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__445__A1 SPB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_404_ _072_ net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__675__A1 DDRA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input28_I io_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__657__A1 _270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_884_ _049_ clknet_3_6__leaf_wb_clk_i PORTB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput23 io_in[12] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput34 io_in[8] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput12 data_in[0] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__662__B _262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__639__A1 _255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__811__A1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__414__I1 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_867_ _032_ clknet_3_2__leaf_wb_clk_i DDRB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_798_ _253_ _376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_721_ PORTA\[1\] _316_ _319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_583_ _201_ _104_ _205_ _209_ _098_ _008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_18_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_652_ _142_ _213_ _267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1 net92 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_49_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I bus_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_704_ DDRB\[5\] _302_ _306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_46_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_566_ _171_ _188_ _189_ _194_ _170_ _006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_635_ net39 _253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_497_ net9 _131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__852__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I DAC_d1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_420_ SPA\[3\] DDRA\[3\] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__875__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_618_ net13 _235_ _240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_549_ _171_ _172_ _175_ _179_ _170_ _004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_42_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__445__A2 DDRB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__898__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_403_ PORTA\[1\] net5 SPA\[1\] _072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__504__I _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_883_ _048_ clknet_3_7__leaf_wb_clk_i PORTB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput13 data_in[1] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput24 io_in[13] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 io_in[9] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input40_I tmr0_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_866_ _031_ clknet_3_0__leaf_wb_clk_i DDRB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_797_ SPA\[5\] _370_ _375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_720_ _270_ _313_ _318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_582_ _206_ _207_ _208_ _209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_9_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__796__A1 net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_651_ _227_ _265_ _266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__720__A1 _270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_849_ _014_ clknet_3_5__leaf_wb_clk_i net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold2 net87 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__787__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__711__A1 DDRB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__702__A1 _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_634_ net17 _235_ _252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_703_ _283_ _292_ _305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_565_ _190_ _191_ _192_ _193_ _194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_496_ net8 _130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__443__S SPB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_617_ net87 _239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_548_ _149_ _176_ _177_ _178_ _179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_39_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_479_ _112_ _113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_14_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_402_ _071_ net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__842__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_38_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_22_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__865__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_882_ _047_ clknet_3_6__leaf_wb_clk_i PORTB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput25 io_in[14] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput14 data_in[2] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput36 pwm0 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__888__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__569__C1 SPA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__408__I0 PORTA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input33_I io_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_865_ _030_ clknet_3_0__leaf_wb_clk_i DDRB\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_796_ net17 _365_ _374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_25_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__903__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_650_ _264_ _265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_581_ SPB\[7\] _154_ _128_ PORTB\[7\] _167_ PORTA\[7\] _208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__583__C _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold3 net89 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_848_ _013_ clknet_3_5__leaf_wb_clk_i net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_779_ _361_ _362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_17_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output64_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_633_ net91 _251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_702_ _181_ _296_ _304_ _254_ _032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_25_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_564_ SPB\[5\] _154_ _123_ net31 _193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_495_ DDRB\[0\] _126_ _128_ PORTB\[0\] _129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__696__A1 _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__448__A1 SPB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__687__A1 _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_616_ _232_ _237_ _238_ _012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_547_ net89 _164_ _103_ _178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_34_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_478_ net6 _112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__678__A1 DDRA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__602__A1 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__669__A1 _248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_401_ _070_ PORTA\[0\] _071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_30_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_881_ _046_ clknet_3_6__leaf_wb_clk_i PORTB\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__814__A1 _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput26 io_in[15] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 data_in[3] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput37 pwm1 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__621__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__408__I1 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__805__A1 _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__531__I _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input26_I io_in[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_864_ _029_ clknet_3_0__leaf_wb_clk_i DDRB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_795_ _372_ _373_ _359_ _056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__855__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_580_ net85 _119_ _143_ DDRA\[7\] _207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__878__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold4 net86 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_847_ _012_ clknet_3_4__leaf_wb_clk_i net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_778_ _360_ _361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__466__A2 _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_632_ _249_ _250_ _238_ _016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_563_ net24 _163_ _164_ net91 _192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_701_ net16 _295_ _304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_494_ _127_ _128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__457__A2 DDRB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__448__A2 DDRB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_615_ _098_ _238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_546_ PORTB\[3\] _128_ _122_ net29 _177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__611__A2 _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_477_ _110_ _111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_400_ SPA\[0\] _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_529_ _093_ _159_ _160_ _081_ _161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_27_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__511__A1 net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__511__B2 DDRA\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_880_ _045_ clknet_3_6__leaf_wb_clk_i PORTB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__578__A1 DDRB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__578__B2 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput27 io_in[1] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput38 pwm2 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput16 data_in[4] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__805__A2 _263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__569__B2 PORTA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input19_I data_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__732__A1 _248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_863_ _028_ clknet_3_0__leaf_wb_clk_i DDRB\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_794_ SPA\[4\] _370_ _373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__723__A1 _242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__542__I _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold5 net88 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_846_ _011_ clknet_3_3__leaf_wb_clk_i net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_777_ _137_ _212_ _360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__475__A3 net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_700_ _301_ _303_ _290_ _031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_631_ net90 _244_ _250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_562_ PORTA\[5\] _167_ _165_ SPA\[5\] _191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__845__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_493_ _112_ _114_ _125_ _127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_1_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_829_ _396_ _397_ _393_ _066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__868__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_46_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_614_ net86 _236_ _237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_545_ net22 _140_ _135_ PORTA\[3\] SPA\[3\] _138_ _176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_39_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_476_ _106_ _109_ _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_54_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__725__I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_459_ _095_ net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__635__I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_528_ _134_ _115_ _130_ _141_ _160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_42_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__511__A2 _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput28 io_in[2] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 rst net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput17 data_in[5] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_862_ _027_ clknet_3_1__leaf_wb_clk_i DDRA\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__420__A1 SPA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_793_ net16 _365_ _372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input31_I io_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold6 net93 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_776_ _357_ _358_ _359_ _051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_845_ _010_ clknet_3_6__leaf_wb_clk_i net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_17_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_29_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_13_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__699__A1 DDRB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_630_ _248_ _231_ _249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_561_ _101_ _149_ _190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_492_ _113_ _121_ _125_ _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_34_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_759_ _275_ _338_ _347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__638__I net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_828_ SPB\[6\] _391_ _397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_613_ _235_ _236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_544_ SPB\[3\] _111_ _173_ DDRB\[3\] _174_ DDRA\[3\] _175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_27_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_475_ _107_ _108_ net8 _109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_33_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__835__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__817__A1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_527_ _134_ _115_ _117_ _141_ _159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_458_ _085_ net21 _095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__858__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput18 data_in[6] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput29 io_in[3] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_43_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_861_ _026_ clknet_3_0__leaf_wb_clk_i DDRA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_792_ _369_ _371_ _359_ _055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_29_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__420__A2 DDRA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input24_I io_in[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold7 net90 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_775_ _322_ _359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_844_ _009_ clknet_3_3__leaf_wb_clk_i net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_17_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_560_ DDRB\[5\] _173_ _174_ DDRA\[5\] _155_ PORTB\[5\] _189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_54_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_491_ net8 _106_ _125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_34_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_30_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__891__CLK clknet_3_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_758_ _086_ _341_ _345_ _346_ _046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_689_ _295_ _296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_827_ _218_ _383_ _396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_612_ _234_ _235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_543_ _142_ _174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__780__A1 _210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_474_ net7 _108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__474__I net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__771__A1 PORTB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__523__A1 SPB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_526_ net45 _158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__753__A1 _270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_457_ _087_ DDRB\[3\] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_10_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput19 data_in[7] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_509_ _142_ _143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_30_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__848__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_860_ _025_ clknet_3_0__leaf_wb_clk_i DDRA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_6_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_791_ SPA\[3\] _370_ _371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__482__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input17_I data_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__410__I0 PORTA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_843_ _008_ clknet_3_4__leaf_wb_clk_i net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output85_I net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold8 net91 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_774_ PORTB\[7\] _351_ _358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__477__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_490_ SPB\[0\] _111_ _120_ net83 _123_ net20 _124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_22_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_826_ _394_ _395_ _393_ _065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_688_ _294_ _295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_757_ _253_ _346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_611_ _132_ _233_ _234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_542_ _126_ _173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_473_ net6 _107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_809_ _110_ _233_ _383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__881__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_456_ _094_ net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__450__A1 _070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_525_ _104_ _148_ _151_ _157_ _147_ _002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__680__A1 _258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__423__A1 SPA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__671__A1 DDRA\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_439_ PORTB\[5\] net2 SPB\[5\] _090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_508_ _141_ _109_ _142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_790_ _360_ _370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__712__B _309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__673__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_3_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__410__I1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_842_ _007_ clknet_3_4__leaf_wb_clk_i net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_773_ _223_ _337_ _357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__838__CLK clknet_3_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__544__C2 DDRA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_756_ net14 _340_ _345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_825_ SPB\[5\] _391_ _395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_687_ _126_ _212_ _294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_610_ _211_ _233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_541_ net46 _172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_472_ net9 _106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_50_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_739_ _255_ _326_ _332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_808_ _082_ _381_ _382_ _147_ _060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_45_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__450__A2 DDRA\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_524_ _152_ _153_ _156_ _157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_455_ _085_ _093_ _094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput90 net102 la_data_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_52_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__423__A2 DDRA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__496__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_438_ _089_ net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_507_ _131_ _141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__871__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__894__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__580__A1 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__571__B2 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__571__A1 PORTB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_772_ _355_ _356_ _349_ _050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_841_ _006_ clknet_3_4__leaf_wb_clk_i net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__562__B2 SPA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__562__A1 PORTA\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__553__B2 _182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__553__A1 _181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__544__A1 SPB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__544__B2 DDRB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_755_ _343_ _344_ _334_ _045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_824_ net17 _384_ _394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_686_ _227_ _292_ _293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__774__A1 PORTB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_540_ _103_ _171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_34_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__765__A1 PORTB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_471_ net43 _105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__517__A1 DDRB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_738_ _330_ _331_ _323_ _041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_669_ _248_ _279_ _280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_807_ _210_ _380_ _382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__756__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__403__S SPA\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_523_ SPB\[1\] _154_ _155_ PORTB\[1\] _156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_output53_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_454_ DDRB\[2\] _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_12_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput80 net80 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput91 net103 la_data_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__729__A1 PORTA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__692__I DDRB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_506_ _107_ _114_ _116_ _106_ _140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_437_ PORTB\[4\] net3 SPB\[4\] _089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_21_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_771_ PORTB\[6\] _351_ _356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_840_ _005_ clknet_3_4__leaf_wb_clk_i net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__861__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__562__A2 _167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__884__CLK clknet_3_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input15_I data_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__808__C _147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output83_I net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_823_ _390_ _392_ _393_ _064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_754_ PORTB\[1\] _341_ _344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_685_ _291_ _292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__628__C _241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_470_ _103_ _104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__517__A2 _126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_806_ _380_ _381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_737_ PORTA\[5\] _328_ _331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_668_ _264_ _279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_599_ net19 _223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_522_ _127_ _155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_453_ _082_ DDRB\[0\] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput70 net70 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__674__A1 _283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput92 net96 la_data_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput81 net81 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__414__S SPA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__665__A1 DDRA\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_436_ _088_ net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_505_ net86 _133_ _136_ PORTA\[0\] SPA\[0\] _138_ _139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_23_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__801__A1 SPA\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_419_ SPA\[1\] DDRA\[1\] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_28_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__647__B _262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_49_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_770_ _218_ _337_ _355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_899_ _064_ clknet_3_3__leaf_wb_clk_i SPB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_31_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_822_ _253_ _393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_753_ _270_ _338_ _343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_684_ _159_ _229_ _291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__851__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_50_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_736_ _283_ _326_ _330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_805_ _110_ _263_ _380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__453__A2 DDRB\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_598_ _099_ _222_ _010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_667_ _276_ _277_ _278_ _023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__874__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__655__B _262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__435__A2 PORTB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_521_ _110_ _154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__897__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_452_ _079_ DDRA\[7\] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_50_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput71 net71 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput93 net101 la_data_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput82 net82 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput60 net60 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_719_ _314_ _317_ _309_ _036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_504_ _137_ _138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_435_ _087_ PORTB\[3\] _088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_3_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input38_I pwm2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_418_ _080_ net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__556__A1 SPB\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_898_ _063_ clknet_3_3__leaf_wb_clk_i SPB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__502__I _135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__710__A1 _258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__777__A1 _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__529__B2 _081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__529__A1 _093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__701__A1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_752_ _339_ _342_ _334_ _044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_821_ SPB\[4\] _391_ _392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__768__A1 PORTB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_683_ _288_ _289_ _290_ _027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__759__A1 _275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_735_ _327_ _329_ _323_ _040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_804_ _079_ _362_ _379_ _346_ _059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_597_ net84 _219_ _221_ _222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_666_ _261_ _278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_520_ net87 _133_ _122_ net27 _144_ _153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__443__I0 PORTB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_451_ _073_ DDRA\[2\] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_35_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput72 net72 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput94 net94 tmr0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput50 net50 data_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput83 net83 irq0 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput61 net61 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_718_ PORTA\[0\] _316_ _317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_649_ _142_ _263_ _264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__841__CLK clknet_3_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__864__CLK clknet_3_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_503_ _107_ _108_ _116_ _106_ _137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_434_ SPB\[3\] _087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__441__S SPB\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__887__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_28_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_417_ _079_ PORTA\[7\] _080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__573__C _098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__902__CLK clknet_3_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_897_ _062_ clknet_3_3__leaf_wb_clk_i SPB\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_751_ PORTB\[0\] _341_ _342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__465__A1 SPA\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_682_ _261_ _290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_820_ _380_ _391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_28_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_44_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__695__A1 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__447__A1 SPB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input13_I data_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__686__A1 _227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_734_ PORTA\[4\] _328_ _329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_803_ _223_ _361_ _379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_665_ DDRA\[3\] _268_ _277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_596_ last_irg6_trigger _220_ _221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__677__A1 _255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I TXD vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_450_ _070_ DDRA\[0\] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_50_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput73 net73 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput95 net95 tmr1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput84 net84 irq6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput51 net51 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput62 net62 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_717_ _315_ _316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__831__A1 SPB\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_648_ _211_ _263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_579_ net93 _164_ _165_ SPA\[7\] _206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_26_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__439__S SPB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_433_ _085_ _086_ net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_502_ _135_ _136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__568__C2 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__521__I _110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_416_ SPA\[7\] _079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_28_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__854__CLK clknet_3_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_42_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_45_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_896_ _061_ clknet_3_3__leaf_wb_clk_i SPB\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__877__CLK clknet_3_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_750_ _340_ _341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__465__A2 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_681_ DDRA\[7\] _281_ _289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_879_ _044_ clknet_3_6__leaf_wb_clk_i PORTB\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__447__A2 DDRB\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_802_ _377_ _378_ _376_ _058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_733_ _315_ _328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_595_ SPB\[0\] net34 _220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_664_ _275_ _265_ _276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__601__A2 _100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__434__I SPB\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput52 net52 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput74 net74 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_716_ _136_ _263_ _315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput85 net85 irq7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput63 net63 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_647_ _259_ _260_ _262_ _019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_578_ DDRB\[7\] _173_ _123_ net33 _204_ _205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
.ends

