* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i
XFILLER_67_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__B1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7963_ _1737_ _3126_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6914_ _2187_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6425__I _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7894_ _4262_ _2334_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A1 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _2068_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5196__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6393__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_3_3__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8515_ _3729_ _3732_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5727_ _4094_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8134__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8446_ _3433_ _1114_ _3426_ _3652_ _3665_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5658_ _4116_ _0840_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ _4189_ _4167_ _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8377_ _3597_ _3598_ _3599_ _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _0993_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7328_ _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8437__A3 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6448__A2 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7259_ _4405_ _2518_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9123__D _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5120__A2 as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5959__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6335__I _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8550__I _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6384__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6136__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7884__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6687__A2 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8833__B1 _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9033__D _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8725__I _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_60_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7939__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4870__A1 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8061__A1 _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _0383_ _0293_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4622__A1 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _4342_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8364__A2 _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _1863_ _1866_ _1877_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_60_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6561_ _1867_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8300_ _2861_ _3511_ _3525_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5512_ _0918_ _0587_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6390__A4 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6492_ _4357_ _4374_ _1808_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8231_ _3422_ _3425_ _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _0771_ _0767_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8162_ _3221_ _3357_ _3390_ _3391_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5350__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ _0548_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7113_ _1789_ _2392_ _2396_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8093_ _2369_ _2666_ _3323_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _4360_ _2335_ _2336_ _0389_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8635__I _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__A1 _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8052__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8995_ _0106_ clknet_leaf_67_wb_clk_i as2650.stack\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6155__I _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _3165_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7877_ _0342_ _4241_ _1252_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5994__I _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8355__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6828_ as2650.r123_2\[2\]\[2\] _2112_ _2141_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6366__A1 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _2073_ _2074_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9118__D _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8429_ _1422_ _3622_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7714__I as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4519__I2 as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7618__A1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7618__B2 _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5234__I _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7094__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8972__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8594__A2 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__A2 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5565__C1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6109__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7857__A1 _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5332__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7085__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ as2650.r123\[3\]\[1\] _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8282__B2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8034__A1 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8585__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7800_ net40 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8780_ _2299_ _3931_ _3936_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5992_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7731_ _0418_ _2969_ _2981_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4943_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7662_ _0405_ _2914_ _1587_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5747__C _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4874_ _4401_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _1910_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6899__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ _2745_ _2845_ _2846_ _2571_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5020__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6544_ _1860_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7848__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7848__B2 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6475_ _1794_ _1786_ _1795_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8214_ _1313_ _1304_ _1296_ _3359_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_133_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5426_ _0571_ _0811_ _0819_ _0834_ _0576_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8145_ _3368_ _3374_ _3260_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5357_ _0629_ _0611_ _0627_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8793__C _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7076__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8076_ _3304_ _3305_ _3306_ _3307_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_87_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5288_ _0663_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5989__I _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__I _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7027_ _2222_ _2316_ _2322_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8995__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6823__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8576__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8978_ _0089_ clknet_leaf_51_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7929_ _3167_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8328__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7709__I _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5011__A1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__A3 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__A4 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8500__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A3 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__I _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5078__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6290__A3 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8224__B _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8319__A2 _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A4 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5139__I _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6750__A1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _4081_ _4183_ _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5553__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _0861_ _1597_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6502__A1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8894__B _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5211_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6191_ net43 _1538_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8255__A1 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ as2650.cycle\[6\] _4260_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8255__B2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5073_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8118__C _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8007__A1 _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8901_ _3185_ _4039_ _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8007__B2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8558__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8832_ _1644_ _3167_ _3171_ _1497_ _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6569__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7230__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _1294_ _1354_ _1358_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8763_ as2650.stack\[4\]\[0\] _3926_ _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7714_ as2650.pc\[9\] _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4926_ _4363_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8694_ _1792_ _3873_ _3878_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7645_ _2840_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _4449_ _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5049__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8730__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8788__C _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7576_ _2809_ _2829_ _2830_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4788_ _4381_ _4229_ _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _0673_ _1842_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7264__I _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8494__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6458_ _1268_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5409_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9177_ _0274_ clknet_leaf_31_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6389_ as2650.psu\[5\] _1501_ _1658_ net28 _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_115_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__A2 _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8128_ _3282_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8797__A2 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8059_ _0398_ _3290_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9173__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8044__B _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__A1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__C _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8182__B1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8721__A2 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5535__A2 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8788__A2 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6518__I _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9041__D _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__I _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__A4 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _1160_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5774__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7793__B _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _4269_ _4053_ _4304_ _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _4204_ _1024_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7430_ _2373_ _2685_ _2686_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8712__A2 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _4225_ _4231_ _4235_ _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6723__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _2346_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4573_ _4134_ _4144_ _4156_ _4166_ _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7084__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _1650_ _0673_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9100_ _0197_ clknet_leaf_37_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8476__A1 _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7279__A2 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7292_ _4434_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9031_ _0142_ clknet_leaf_20_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6243_ _1578_ _1420_ _1584_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8491__A4 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _0317_ _4338_ _1521_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__8228__B2 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5125_ _0531_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6428__I _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7451__A2 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5056_ _4086_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7968__B _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5462__A1 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7687__C _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6006__A3 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8815_ _3250_ _3303_ _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__A1 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8746_ _3901_ _2141_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6962__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ as2650.stack\[2\]\[7\] _1341_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4909_ as2650.cycle\[0\] _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5889_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8677_ _2291_ _3865_ _3867_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8703__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7628_ _1327_ _1140_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7559_ _1587_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5507__I _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8219__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7690__A2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6338__I _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__I _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7442__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_7__f_wb_clk_i clknet_0_wb_clk_i clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9069__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__B1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8502__B _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5508__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9036__D _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7632__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6248__I _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5152__I _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8891__C _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4991__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7984__A3 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6930_ _4081_ _1811_ _2239_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6861_ _2116_ _2139_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7197__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__I as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8394__B1 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8600_ _3687_ _1177_ _3810_ _3811_ _2814_ _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5812_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6792_ _0875_ _2098_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6944__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5747__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__I0 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8531_ _3736_ _3747_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5743_ _1139_ _1026_ _1146_ _0879_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8462_ _3487_ _1128_ _3551_ _3670_ _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5674_ _4172_ _4175_ _4133_ _0942_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7413_ _2665_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _4212_ _4214_ _4216_ _4218_ _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8393_ _2374_ _3590_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6172__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__I _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _2592_ _2551_ _2600_ _2602_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8449__A1 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _4149_ _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7970__C _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ _2527_ _0321_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _4069_ _4074_ _4080_ _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7121__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6226_ _0699_ _0708_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9014_ _0125_ clknet_leaf_34_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7672__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4486__A2 _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6157_ _4440_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5108_ _4356_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7424__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8621__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _1450_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5435__A1 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _0413_ _0300_ _0415_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A3 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__B _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6935__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8729_ _3902_ _3903_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8929__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6163__A2 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5237__I as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput20 net20 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_108_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput31 net31 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8860__A1 _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A1 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6068__I _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7966__A3 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__S _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6926__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6387__C1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7627__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8679__A1 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7351__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A2 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ as2650.addr_buff\[6\] _0653_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4986__I _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ _2352_ _4346_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _1370_ _1386_ _1388_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8603__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7962_ _3198_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5610__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6913_ _2173_ _2195_ _2196_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_70_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7893_ _4423_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6844_ _4099_ _1864_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6775_ _2071_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6441__I _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8514_ _0698_ _3731_ _2482_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5726_ _0743_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8445_ _3194_ _3659_ _3664_ _0435_ _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5657_ as2650.holding_reg\[5\] _0595_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4608_ _4173_ _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8376_ _2497_ _0908_ _3551_ _3582_ _3495_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5588_ _0987_ _0991_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4546__I3 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7327_ _2585_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4539_ _4129_ _4132_ _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8842__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7258_ _2493_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A1 _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__B _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _1529_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7189_ _2458_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7221__B _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A1 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__B1 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6384__A2 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6136__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__B1 _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7884__A2 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__I3 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7636__A2 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8833__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8833__B2 _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A3 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A2 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8061__A2 _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6072__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A2 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _0318_ _0293_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7947__I0 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__B1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7572__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6560_ _1870_ _1873_ _1876_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8897__B as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5511_ _4128_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6491_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8230_ _2782_ _3457_ _3313_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5442_ _0848_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7875__A2 _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__I3 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8161_ _3219_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5373_ _4215_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7092__I _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ as2650.stack\[4\]\[9\] _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8092_ _3027_ _3322_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8824__A1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7043_ _1245_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7820__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8588__B1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4861__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8052__A2 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8994_ _0105_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__A1 as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7945_ _0970_ _3174_ _3184_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7876_ _3120_ _3102_ _3121_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_35_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _2037_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7563__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6366__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7267__I _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _4076_ _1902_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ _0831_ _1111_ _1112_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7315__A1 _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6689_ _4106_ _2005_ _1975_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8428_ _0333_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7866__A2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4519__I3 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8359_ _3581_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__B _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8815__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8291__A2 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8579__B1 _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5250__I _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__B1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6109__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__B1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7857__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7126__B _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9044__D _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8806__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6293__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ _2678_ _2977_ _2980_ _2808_ _0417_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _4397_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7661_ _2881_ _2913_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4873_ _4370_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7545__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7087__I _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8742__B1 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6612_ _0776_ _1922_ _1923_ _0876_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7592_ _1673_ _2568_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6899__A3 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6543_ as2650.r123\[0\]\[4\] as2650.r123_2\[0\]\[4\] _4088_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7848__A2 _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ as2650.stack\[6\]\[11\] _1790_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5859__A1 _4439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8213_ _3276_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5425_ _0743_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5335__I _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8144_ _0376_ _3369_ _3373_ _3128_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5356_ _0764_ _0755_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8646__I _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8075_ as2650.stack\[1\]\[1\] _3242_ _3254_ as2650.stack\[0\]\[1\] _0722_ _3307_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_47_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6284__A1 _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7026_ as2650.r123_2\[1\]\[5\] _2304_ _2320_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5070__I _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6036__A1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8977_ _0088_ clknet_leaf_51_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7784__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7784__B2 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ _3170_ _1676_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _2487_ _3102_ _3104_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__7536__A1 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6115__B _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5011__A2 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6511__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__I _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5078__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8016__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6027__A1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7775__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8505__B _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__C _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7527__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__B2 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__A2 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6502__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0614_ _4230_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4513__A1 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6190_ _1540_ _1533_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4994__I _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5141_ _0549_ _4310_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8255__A2 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7370__I _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _4079_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8900_ _3184_ _4037_ as2650.psu\[3\] _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8007__A2 _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6018__A1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8831_ _3982_ _3939_ _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7766__A1 as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8762_ _3924_ _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5974_ as2650.stack\[1\]\[2\] _1355_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7713_ _2787_ _2963_ _2964_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8693_ as2650.stack\[5\]\[10\] _3876_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8715__B1 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7644_ _2879_ _2729_ _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4856_ _4419_ _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7575_ _0350_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4787_ _4302_ _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6526_ _0674_ _1811_ _1838_ _1841_ _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8494__A2 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6457_ _1385_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8962__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5408_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9176_ _0273_ clknet_leaf_31_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6388_ _1723_ _1021_ _1724_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ _1298_ _3356_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7049__A3 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _0694_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6257__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8058_ _1287_ _2536_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _1927_ _2308_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_6__f_wb_clk_i clknet_0_wb_clk_i clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7757__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5232__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output12_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7509__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7455__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8485__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5299__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6496__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8286__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7190__I _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7996__A1 _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5223__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _4302_ _4303_ _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8173__A1 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5690_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__B _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4989__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _4232_ _4225_ _4234_ _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6723__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7920__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7360_ _2613_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4572_ _4157_ _4158_ _4165_ _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6311_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7291_ _2550_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9030_ _0141_ clknet_leaf_20_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6242_ as2650.stack\[3\]\[12\] _1580_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ _4430_ _0325_ _4335_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5613__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _0532_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5055_ _0472_ _0473_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_73_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7739__A1 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8145__B _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6444__I _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8814_ _3958_ _3966_ _3967_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7984__B _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8745_ _0901_ _3911_ _3912_ as2650.r123\[2\]\[2\] _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5957_ _1325_ _1340_ _1344_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4908_ _4243_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8676_ as2650.stack\[6\]\[4\] _3866_ _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8164__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ _0753_ _1288_ _1281_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7627_ _2529_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4839_ _4431_ _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7911__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6714__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4725__A1 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _2795_ _2807_ _2812_ _2607_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7489_ _2568_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__A1 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9140__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7224__B _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8219__A2 _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9159_ _0256_ clknet_leaf_6_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5523__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6354__I _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6402__A1 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8502__C _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7902__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__A2 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7185__I _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6957__C _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5692__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6641__A1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__B _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6860_ _2172_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8394__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7197__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8394__B2 _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5811_ net3 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _0877_ _2042_ _1835_ _2105_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6944__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8530_ _1541_ _1615_ _3744_ _3746_ _3727_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5742_ _1143_ _1024_ _1145_ _0685_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8146__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8461_ _0395_ _3677_ _3678_ _3679_ _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7095__I _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5673_ _0583_ _1059_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8697__A2 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7412_ _1764_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4707__A1 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9163__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4209_ _4217_ _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8392_ _3607_ _3613_ _3232_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7343_ _2601_ _2365_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5380__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ as2650.r0\[1\] _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7274_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4486_ _4076_ _4079_ _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7121__A2 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9013_ _0124_ clknet_leaf_35_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6225_ _1554_ _1570_ _1571_ _1568_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6439__I _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__I _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _4300_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6883__B _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _4064_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7424__A3 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6087_ as2650.r123_2\[3\]\[0\] _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8621__A2 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6632__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5435__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5038_ _0339_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input11_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8385__A1 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ as2650.stack\[5\]\[4\] _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8728_ _1108_ _3893_ _3890_ as2650.r123\[1\]\[5\] _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8137__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8322__C _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8659_ as2650.stack\[7\]\[13\] _3847_ _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8688__A2 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6163__A3 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5371__A1 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7112__A2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5253__I _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5674__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8073__B1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8612__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__A2 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__B1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6387__C2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9186__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8232__C _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5428__I as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7351__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__A1 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6010_ as2650.stack\[1\]\[8\] _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8603__A2 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5417__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7961_ _3197_ as2650.holding_reg\[6\] _3186_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6912_ _2179_ _2194_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7892_ _2500_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8367__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _0988_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6774_ _2075_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8513_ _3730_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _0820_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5338__I as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8444_ _2472_ _3654_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5656_ _4115_ _0540_ _1060_ _4376_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5353__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _4171_ _4180_ _4200_ _4173_ _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8375_ _3339_ _3582_ _3555_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7553__I _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7326_ _2584_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4538_ _4071_ _4130_ _4131_ _4068_ _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_89_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__A1 as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7257_ _0731_ _2509_ _2516_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4469_ _4062_ _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5073__I _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8842__A2 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _1303_ _1555_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5900__I0 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7188_ _2457_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9059__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6139_ _4298_ _4390_ _4369_ _0631_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_100_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6081__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8358__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__A1 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__B2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7581__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7463__I _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7097__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__A1 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8349__A1 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7947__I1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5583__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _0602_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6490_ _4082_ _0516_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _0842_ _0847_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7875__A3 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8160_ _3377_ _3389_ _2731_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5372_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _2390_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8091_ _3319_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8824__A2 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6835__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7042_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8588__A1 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8588__B2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8993_ _0104_ clknet_leaf_59_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A1 _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7944_ _4362_ _1680_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7976__C _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7875_ _4267_ _4275_ _2518_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7012__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _2114_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7563__A2 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8760__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _2022_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5574__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ as2650.stack\[5\]\[13\] _0824_ _0827_ as2650.stack\[4\]\[13\] _0825_ _1113_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_136_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _1906_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7315__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8600__C _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8427_ _3624_ _3646_ _3647_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5639_ as2650.stack\[7\]\[12\] _1043_ _1044_ as2650.stack\[6\]\[12\] _1045_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7866__A3 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__I _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8358_ _1400_ _3580_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7309_ _1708_ _0650_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8289_ _4262_ _4435_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8815__A2 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8579__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A1 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7251__B2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7458__I _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6362__I _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__B1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8751__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6109__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8503__A1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8510__C _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7193__I _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7126__C _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8806__A2 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7490__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6537__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6293__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _0707_ _1348_ _1366_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _4365_ _0363_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7660_ _2854_ _2858_ _2882_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4872_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7545__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8742__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6611_ _1905_ _1926_ _1927_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5556__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7591_ _2841_ _2844_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6542_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _1413_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5616__I _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8212_ _0437_ _0679_ _3435_ _3439_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5859__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _0820_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9192_ _0289_ clknet_leaf_45_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8143_ _1679_ _3292_ _3370_ as2650.addr_buff\[3\] _3372_ _0398_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_5355_ as2650.holding_reg\[1\] _0585_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6808__A1 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8074_ as2650.stack\[3\]\[1\] _3302_ _3303_ as2650.stack\[2\]\[1\] _3306_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5286_ _0580_ _0638_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7481__A1 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7025_ _1854_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6284__A2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_wb_clk_i clknet_0_wb_clk_i clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7233__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8976_ _0087_ clknet_leaf_51_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7784__A2 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7927_ _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7858_ _2555_ _0420_ _1482_ _2344_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_51_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7536__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8733__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _2082_ _2086_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5547__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7789_ _3009_ _2786_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6910__I _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7942__S _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8058__B _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6357__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5078__A3 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7897__B _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_79_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7775__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5786__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7188__I _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__B _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4541__S _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__A2 _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__I _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4513__A2 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _0515_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5071_ _0481_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__A1 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8830_ _3176_ _1644_ _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7766__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8761_ _3924_ _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5973_ _1290_ _1354_ _1357_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7098__I _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7712_ _2931_ _2829_ _2830_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4515__I _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _4343_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8692_ _1789_ _3873_ _3877_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8715__B2 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7643_ _4443_ _2895_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5529__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _4447_ _4448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7574_ _2524_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4786_ _4374_ _4379_ _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6525_ _4449_ _0546_ _1809_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_101_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _1434_ _1772_ _1780_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _0814_ _0815_ _0560_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9175_ _0272_ clknet_leaf_31_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7561__I _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6387_ _0708_ _1712_ _1718_ as2650.psu\[2\] as2650.psu\[7\] _1214_ _1725_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_8126_ as2650.pc\[2\] _2582_ _1274_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_86_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5338_ as2650.r123\[0\]\[1\] _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6177__I _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8057_ _2263_ _2590_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _4045_ _4344_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _1897_ _2307_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8606__B _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7206__A1 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5768__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8959_ _0070_ clknet_leaf_66_wb_clk_i as2650.r123_2\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7937__S _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__A3 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__A2 _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8706__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8182__A2 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7693__A1 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6496__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7445__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7996__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4536__S _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__A2 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6708__B1 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8173__A2 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4640_ _4053_ _4233_ _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_124_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7920__A2 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4734__A2 _4327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _4164_ _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6310_ _0666_ _0448_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7290_ _4430_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6241_ _1577_ _1414_ _1583_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7381__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _1521_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5123_ as2650.addr_buff\[5\] _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6239__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _4381_ _4234_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6725__I _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7739__A2 _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8813_ _2280_ _3958_ _0351_ _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8744_ _3913_ _3914_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ as2650.stack\[2\]\[6\] _1341_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8675_ _3858_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5887_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7626_ as2650.pc\[7\] _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4838_ _4430_ _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6175__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7557_ _2808_ _2811_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4725__A2 _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5076__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _4362_ _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _0543_ _1260_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7488_ _0639_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7675__A1 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6478__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6439_ _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7291__I _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__A1 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9158_ _0255_ clknet_leaf_73_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8109_ _1489_ _3327_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9089_ _0186_ clknet_leaf_17_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6650__A2 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5695__B _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7466__I _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8155__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7902__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7666__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7130__A3 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A2 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7418__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_23_wb_clk_i clknet_opt_4_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4493__C _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8952__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5810_ _1212_ _0782_ _0612_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_63_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6790_ _0674_ _2045_ _2099_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6944__A3 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _1144_ _0683_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8146__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6280__I _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8460_ _2382_ _3463_ _3235_ _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5672_ _1004_ _1068_ _1072_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6157__A1 _4440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7411_ _2666_ _2632_ _2667_ _2668_ _1259_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _4194_ _4210_ _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8391_ _3473_ _3609_ _3611_ _3162_ _3612_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4707__A2 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7342_ _2554_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _4147_ _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5380__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7657__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7273_ _2531_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4485_ _4078_ _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9012_ _0123_ clknet_leaf_34_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6224_ net22 _1559_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A1 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6155_ _4342_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8082__A1 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _4309_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6086_ _1331_ _1444_ _1449_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _0436_ _0439_ _0441_ _0444_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6632__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5499__C _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8385__A2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6396__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6988_ _2281_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8727_ _3901_ _2320_ _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__A2 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _1243_ _0705_ _1270_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8137__A2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4703__I _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8658_ _1796_ _3849_ _3855_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7896__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _4447_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8589_ _2144_ _1696_ _0520_ _1668_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5371__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5534__I _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A1 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6387__B2 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4613__I _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6139__A1 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7887__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7639__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__A1 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8064__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7811__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6275__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7960_ _1122_ _3174_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4625__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6911_ _2190_ _2193_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7891_ _2503_ _3122_ _3125_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_78_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _2003_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9130__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8423__C _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6773_ _2078_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5050__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ _1124_ _1125_ _1126_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8512_ _3726_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7878__A1 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_4_0_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8443_ _3339_ _3658_ _3662_ _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5655_ _4106_ _0587_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4606_ _4126_ _4195_ _4199_ _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8374_ _3188_ _3585_ _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6550__A1 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ _0987_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7325_ net3 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4537_ as2650.r123\[1\]\[3\] as2650.r123\[0\]\[3\] as2650.r123_2\[1\]\[3\] as2650.r123_2\[0\]\[3\]
+ _4058_ _4110_ _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7256_ _1279_ _2515_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6302__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__A2 as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _4061_ _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _1099_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8665__I _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7187_ _1366_ _2456_ _1367_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5900__I1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8055__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6138_ _4374_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ as2650.stack\[0\]\[0\] _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4616__A1 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8614__B _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8333__C _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8987__D _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8530__A2 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5264__I _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8294__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7097__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9003__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__A2 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9153__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7919__I _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5032__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6780__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _0842_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6532__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ _4413_ _0526_ _0536_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5174__I as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7110_ _1781_ _2392_ _2394_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8285__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8090_ _3283_ _3284_ _3320_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7041_ _4447_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8037__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8588__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_4__f_wb_clk_i clknet_0_wb_clk_i clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8992_ _0103_ clknet_leaf_59_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout54_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7260__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _3183_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5271__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6733__I _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5777__C _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _0434_ _2518_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7012__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _2116_ _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5023__A1 _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8760__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ _4138_ _1973_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ as2650.stack\[7\]\[13\] _1043_ _1044_ as2650.stack\[6\]\[13\] _1112_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6687_ _0662_ _2003_ _1971_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8426_ _0469_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5638_ _0717_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7866__A4 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8357_ as2650.pc\[9\] _1378_ _3530_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5569_ _0906_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7308_ _0641_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8288_ _1328_ _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8609__B _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7239_ _2497_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__I _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9176__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8028__A1 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8344__B _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8751__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__A1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7474__I _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5317__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8267__A1 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7490__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4940_ _0364_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5005__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5169__I _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8742__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _0776_ _0589_ _1922_ _1898_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_127_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7590_ _2842_ _2804_ _2843_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5556__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9049__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4801__I _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6472_ _1792_ _1786_ _1793_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6505__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6221__C _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8211_ _3424_ _3436_ _3438_ _2330_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5423_ _0823_ _0826_ _0830_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5859__A3 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9191_ _0288_ clknet_leaf_45_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8258__A1 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8142_ _1297_ _1216_ _3371_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5354_ _4148_ _4154_ _4394_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6808__A2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8073_ as2650.stack\[5\]\[1\] _2456_ _3254_ as2650.stack\[4\]\[1\] _0906_ _3305_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_99_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5285_ _0644_ _0651_ _0693_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4819__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7024_ _1937_ _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7481__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7233__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8975_ _0086_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7559__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__I _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7926_ _3168_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5795__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7857_ _4337_ _0330_ _3103_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_90_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8733__A2 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6808_ _4100_ _1915_ _2087_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6744__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7788_ _0350_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7508__B _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _0753_ _2042_ _2043_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7294__I _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5807__I _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8497__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8409_ _3401_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8249__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5542__I _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5078__A4 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A2 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8421__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5786__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__B1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5717__I _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7160__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7932__I _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _4391_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__A2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8412__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6283__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8760_ _2280_ _0715_ _1270_ _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ as2650.stack\[1\]\[1\] _1355_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7711_ _1381_ _2880_ _2962_ _0340_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4923_ _0333_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8691_ as2650.stack\[5\]\[9\] _3876_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8715__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7642_ _2879_ _0377_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4854_ _4274_ _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5529__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7573_ _2789_ _2530_ _2815_ _0458_ _2827_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_105_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4785_ _4378_ _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4531__I _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _1839_ _1840_ _1810_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6455_ as2650.stack\[0\]\[14\] _1770_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5406_ _0488_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6386_ _0699_ _1708_ _1709_ as2650.psu\[3\] _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_9174_ _0271_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8125_ _3353_ _3355_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5337_ _0514_ _0578_ _0746_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6458__I _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8056_ _2353_ _3286_ _3287_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5268_ _4322_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5465__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7007_ _0778_ _1923_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ as2650.psl\[3\] _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7206__A2 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8403__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6193__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8958_ _0069_ clknet_leaf_61_wb_clk_i as2650.r123_2\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7909_ _0315_ _2495_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8889_ _3178_ _4030_ _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8706__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7390__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7953__S _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7693__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8069__B _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5272__I _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7445__A2 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7701__B _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6956__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__A3 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8532__B _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7927__I _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _4163_ _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5931__A2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7133__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ as2650.stack\[3\]\[11\] _1580_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5695__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6171_ _1524_ _4445_ _0381_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5122_ as2650.addr_buff\[6\] _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8633__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7611__B _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _4396_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8812_ _3964_ _3965_ _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8743_ _3901_ _2094_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _1317_ _1340_ _1343_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6741__I _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4906_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8674_ _3858_ _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5886_ as2650.pc\[1\] _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7625_ _0335_ _2878_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4837_ _4411_ _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7556_ _2809_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_105_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5922__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ _4361_ _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6507_ _4284_ _0419_ _1803_ _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7487_ _0406_ _2698_ _2742_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4699_ _4238_ _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8872__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6438_ _0700_ _1348_ _1351_ _1367_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__4489__A2 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6188__I _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9157_ _0254_ clknet_leaf_3_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _1702_ _1703_ _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_121_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8108_ _1474_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9088_ _0185_ clknet_leaf_16_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5438__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8039_ _3219_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4661__A2 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6651__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7115__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8863__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5677__A1 _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A3 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7418__A2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8615__A1 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5429__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6929__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5601__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__B2 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5740_ _4104_ _4187_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7354__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5177__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5671_ _0931_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6157__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7410_ _2630_ _0461_ _2355_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4622_ _4158_ _4215_ _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8390_ _3436_ _3603_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7341_ _2552_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4553_ _4146_ _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5905__I _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7272_ _0813_ _4439_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4484_ _4077_ _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8854__A1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9011_ _0122_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6223_ _1240_ _1555_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A2 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _1458_ _1487_ _1506_ _1508_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8606__A1 _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ as2650.cycle\[0\] as2650.cycle\[8\] _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ as2650.stack\[0\]\[7\] _1445_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5640__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _4371_ _0450_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__B2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6987_ _2281_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8726_ _3900_ _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _1302_ _1331_ _1332_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4946__A3 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__C _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8657_ as2650.stack\[7\]\[12\] _3851_ _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5087__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__A1 _4437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5869_ _1243_ _0719_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8900__B as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6148__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7608_ _2832_ _0461_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7896__A2 _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8588_ _1864_ _0502_ _3432_ _0732_ _1700_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7539_ _2790_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5371__A3 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8845__A1 _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput12 net12 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5659__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 net23 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput45 net45 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8073__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__A1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_0__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__B1 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7584__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6387__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A3 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6314__C _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7336__A1 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6139__A2 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7887__A2 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9082__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7639__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8836__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4873__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_3__f_wb_clk_i clknet_0_wb_clk_i clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8064__A2 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7811__A2 _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__A2 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8771__I _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7890_ _3101_ _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _2118_ _2138_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _2012_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8511_ _3694_ _3728_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ as2650.stack\[3\]\[14\] _1043_ _1044_ as2650.stack\[2\]\[14\] _0973_ _1127_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8442_ _3512_ _3659_ _3661_ _3278_ _3033_ _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7878__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5654_ _1055_ _4379_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _4129_ _4132_ _4137_ _4142_ _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8373_ _3593_ _3595_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5585_ as2650.holding_reg\[4\] _0917_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7324_ _2529_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4561__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4536_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _4110_ _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _4298_ _0491_ _0486_ _0501_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ as2650.psl\[4\] _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6302__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _1532_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4695__B _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7186_ _2455_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6466__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8055__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _1088_ _4361_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5370__I _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _1437_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__A2 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5019_ _0437_ _0394_ _0438_ _0300_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8614__C _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__I _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8709_ _3885_ _1924_ _3888_ as2650.r123\[1\]\[0\] _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7318__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7869__A2 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5545__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7961__S _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8818__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8294__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4607__A2 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5280__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_4_0_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_opt_4_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7557__A1 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5568__B1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5568__C2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__A2 _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__A2 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8809__A1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _0545_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8285__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7040_ _2331_ _1764_ _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8037__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8991_ _0102_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__A2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7942_ _3182_ as2650.holding_reg\[2\] _3166_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7873_ net50 _3116_ _3119_ _2629_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8745__B1 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4534__I _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _2118_ _2138_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__A2 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _2017_ _2069_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ as2650.stack\[3\]\[13\] _0821_ _0718_ as2650.stack\[2\]\[13\] _1110_ _1111_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_52_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _1973_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8425_ _3273_ _3627_ _3645_ _3622_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5637_ _0714_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6523__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8356_ _1390_ _3499_ _3579_ _0349_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5568_ as2650.stack\[5\]\[11\] _0704_ _0710_ as2650.stack\[4\]\[11\] as2650.stack\[7\]\[11\]
+ _0713_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7307_ _2329_ _2565_ _2566_ _0419_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4519_ as2650.r123\[1\]\[5\] as2650.r123\[0\]\[5\] as2650.r123_2\[1\]\[5\] as2650.r123_2\[0\]\[5\]
+ _4059_ _4063_ _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8287_ _1320_ _3442_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5499_ as2650.stack\[1\]\[10\] _0824_ _0827_ as2650.stack\[0\]\[10\] _0906_ _0907_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_137_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _1247_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__B _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8028__A2 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7169_ _1114_ _2428_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6129__C _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7787__A1 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__A1 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__A2 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8751__A3 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5275__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__B2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5722__B1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8267__A2 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6278__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8519__C _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5325__I0 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7778__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _4226_ _4420_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5005__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7950__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8988__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6540_ as2650.r123\[0\]\[5\] as2650.r123_2\[0\]\[5\] as2650.psl\[4\] _1857_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6471_ as2650.stack\[6\]\[10\] _1790_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7702__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _1501_ _4448_ _3437_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5422_ _0722_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9190_ _0287_ clknet_leaf_43_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8141_ _2263_ _2717_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5353_ _0758_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6269__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6808__A3 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8072_ as2650.stack\[7\]\[1\] _3302_ _3303_ as2650.stack\[6\]\[1\] _3304_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5284_ _0567_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4819__A2 _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7023_ _1920_ _1935_ _1936_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_87_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8974_ _0085_ clknet_leaf_16_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _4047_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8718__B1 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7856_ _4334_ _2492_ _2494_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _0918_ _2003_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7575__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7787_ _3000_ _2880_ _3036_ _2996_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4999_ as2650.cycle\[2\] _0296_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6744__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _2044_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8497__A2 _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6669_ _4149_ _1858_ _4091_ _4159_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8408_ _2378_ _3628_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4507__A1 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__B1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9143__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8249__A2 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8339_ _1389_ _3533_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5180__A1 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5483__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8421__A2 _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__A1 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__B2 as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4746__A1 _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__B _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_17_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6499__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8660__A2 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6671__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8412__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__B2 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _1284_ _1354_ _1356_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9016__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7710_ _2935_ _2944_ _2960_ _2961_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4985__A1 _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4922_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8690_ _3871_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8176__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7641_ _2600_ _2890_ _2893_ _2331_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4853_ _4364_ _4445_ _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5908__I _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__I _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _2816_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4784_ _4377_ _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _0680_ _1808_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8479__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _1427_ _1772_ _1779_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7344__B _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5162__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9173_ _0270_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ as2650.psu\[4\] _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8159__C _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8124_ _2664_ _3269_ _3354_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _0579_ _0697_ _0735_ _0744_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8100__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8055_ _0787_ _2334_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8651__A2 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5267_ _0370_ _4326_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7006_ _2303_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6662__A1 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5198_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8957_ _0068_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7908_ _1588_ _3152_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4976__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8167__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8888_ _3976_ _4028_ as2650.psl\[1\] _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7839_ _3022_ _3080_ _3082_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7914__A1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7390__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5039__B _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5153__A1 _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8642__A2 _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6653__B2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6405__A1 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7602__B1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8813__B _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6420__A4 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9189__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8158__A1 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6169__B1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5392__A1 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7133__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5144__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8881__A2 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__I _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__A1 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__A2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6170_ _4359_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5121_ _0529_ _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5447__A2 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5052_ _4085_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__I _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8811_ _3258_ _0723_ _3960_ _0424_ _3965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8742_ _0811_ _3911_ _3912_ as2650.r123\[2\]\[1\] _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5954_ as2650.stack\[2\]\[5\] _1341_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__C _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7339__B _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4905_ _0322_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8673_ _2289_ _3859_ _3864_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__I _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5885_ _1272_ _1284_ _1286_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7624_ _2832_ _2581_ _2877_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4836_ _4424_ _4428_ _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6175__A3 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7555_ net33 _2741_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4767_ _4360_ _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ as2650.cycle\[9\] _4281_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7486_ _2740_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8321__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4698_ _4259_ _4291_ _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5135__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6437_ _1768_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5373__I _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8872__A2 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9156_ _0253_ clknet_leaf_6_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6368_ _1679_ _4207_ _4209_ _0786_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8107_ _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ as2650.stack\[3\]\[8\] _0715_ _0719_ as2650.stack\[2\]\[8\] _0728_ _0729_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_62_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9087_ _0184_ clknet_leaf_23_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6299_ _4359_ _0448_ _0290_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _3267_ _3270_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4717__I _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8388__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6938__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7060__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7964__S _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4452__I _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7115__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5677__A2 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2__f_wb_clk_i clknet_0_wb_clk_i clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6626__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8527__C _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7003__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8379__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8543__B _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7051__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6842__I _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8262__C _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _1066_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8551__A1 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5365__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _4165_ _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _2592_ _2540_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7606__C _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4552_ _4067_ _4145_ _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8303__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5117__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7271_ _0376_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ _4066_ as2650.ins_reg\[1\] _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9010_ _0121_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6865__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _1139_ _1556_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6153_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8606__A2 _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ as2650.r123\[0\]\[0\] _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6084_ _1325_ _1444_ _1448_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _0299_ _0453_ _0446_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8009__I _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _1308_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7593__A2 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8790__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8725_ _0741_ _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5937_ as2650.stack\[3\]\[7\] _1310_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8656_ _1794_ _3848_ _3854_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5868_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7345__A2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8542__A1 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7607_ _4440_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4819_ as2650.cycle\[3\] _4411_ _4412_ _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5356__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8587_ as2650.psl\[5\] _3698_ _1460_ _3799_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7896__A3 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _1161_ _1176_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7538_ _2791_ _2792_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7516__C _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5108__A1 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6199__I _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7469_ _2722_ _2697_ _2725_ _0440_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8845__A2 _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 net13 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5659__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput46 net46 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9139_ _0236_ clknet_leaf_44_wb_clk_i as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6927__I _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5831__I _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6608__A1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7251__C _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6084__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8363__B _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__A1 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7033__B2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8082__C _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8781__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7336__A2 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8810__C _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7887__A3 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4910__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8836__A2 _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8049__B1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8257__C _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7272__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6075__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__A3 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5822__A2 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6840_ _2121_ _2137_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5035__B1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2082_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8510_ _1534_ _1615_ _3707_ _3708_ _3727_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_52_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5722_ as2650.stack\[1\]\[14\] _0705_ _0711_ as2650.stack\[0\]\[14\] _1126_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8524__A1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8441_ _3650_ _3660_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5653_ _1056_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7878__A3 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _4189_ _4197_ _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8372_ _3537_ _3582_ _3594_ _3278_ _3033_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5584_ _4125_ _0541_ _0989_ _4377_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ as2650.pc\[1\] _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4535_ _4128_ _4078_ _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4561__A2 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6838__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7254_ _2512_ _2513_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4466_ _4059_ _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6205_ _1532_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__I as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4695__C _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _1489_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7263__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5018_ _4242_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7578__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8763__A1 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _1831_ _2272_ _2277_ _2278_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8708_ _3887_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8639_ _2295_ _3840_ _3843_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__I _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5047__B _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8279__B1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8818__A2 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6829__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__I _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9180__D _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__A1 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8093__B _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7488__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4905__I _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8203__B1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7557__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8821__B _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8506__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7309__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4791__A2 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8809__A2 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6296__A2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__I0 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5471__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9090__D _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7245__A1 _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8990_ _0101_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7941_ _3180_ _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4815__I _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7872_ _3116_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7548__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8745__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _2121_ _2137_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5559__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _2019_ _2031_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5705_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ _2000_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4550__I _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8424_ _3643_ _3644_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5636_ as2650.stack\[1\]\[12\] _0725_ _0822_ as2650.stack\[2\]\[12\] _1041_ _1042_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_104_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8355_ _3422_ _3562_ _3578_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5567_ as2650.stack\[3\]\[11\] _0715_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5731__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7306_ _0326_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4518_ _4072_ _4111_ _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8286_ _3281_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7237_ _1512_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5495__B1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ _2441_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7236__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7099_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9072__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8736__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7257__B _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4460__I as2650.alu_op\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__A2 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A1 as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__B2 as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5492__S _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7475__A1 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6278__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7475__B2 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5325__I1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5291__I as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8816__B _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7227__A1 _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7778__A2 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__A2 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8727__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7946__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5005__A3 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8270__C _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7950__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6470_ _1403_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ as2650.stack\[0\]\[9\] _0827_ _0718_ as2650.stack\[2\]\[9\] _0829_ _0830_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ _3293_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5352_ _0758_ _0760_ _0621_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8071_ _1573_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5283_ _0652_ _0660_ _0691_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ _2209_ _2316_ _2318_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9095__CLK clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__B _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7218__A1 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8445__C _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8973_ _0084_ clknet_leaf_16_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4545__I _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8017__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7924_ _0663_ _1463_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8718__B2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7855_ _1626_ _1247_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8932__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6806_ _2075_ _2089_ _2120_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7786_ _3013_ _3021_ _3035_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4998_ _0413_ _0418_ _0420_ _4432_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7941__A2 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6737_ _0782_ _2045_ _2052_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5376__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6668_ as2650.r0\[1\] _4089_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7805__B _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8407_ as2650.addr_buff\[2\] as2650.addr_buff\[3\] _3589_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8687__I _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5619_ _4198_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4507__A2 _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ _0588_ _1915_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8338_ _3561_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7457__A1 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8269_ _3487_ _3493_ _3494_ _3495_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4455__I _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8185__A2 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4746__A2 _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5943__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__A3 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7696__A1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6499__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__A2 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7006__I _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6120__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6671__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8412__A3 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8955__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7620__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ as2650.stack\[1\]\[0\] _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ as2650.cycle\[8\] _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4985__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7640_ net54 _2821_ _2891_ _2892_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4852_ _4323_ _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5529__A4 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7571_ _1314_ _2534_ _2825_ _2729_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4737__A2 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4783_ _4376_ _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5934__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _4158_ _4215_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8479__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6453_ as2650.stack\[0\]\[13\] _1770_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5404_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9172_ _0269_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5162__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6384_ _1465_ _1467_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7439__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8123_ _1686_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5335_ _0576_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8054_ _3283_ _3284_ _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6111__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7005_ _1852_ _2302_ _2305_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _0594_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7611__A1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8956_ _0067_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _0299_ _2492_ _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4976__A2 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8191__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8887_ _4032_ _4033_ _3647_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8167__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6178__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7838_ _4410_ _3085_ _2943_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7769_ _3017_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7678__A1 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7678__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6350__A1 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4900__A2 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_1__f_wb_clk_i clknet_0_wb_clk_i clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_79_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7850__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8978__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__A1 _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7602__A1 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6405__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8158__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4913__I as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6169__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7905__A2 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5392__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7669__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8866__B1 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8120__I _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5120_ _4386_ as2650.cycle\[8\] _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__A1 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6644__A2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5051_ _0428_ _4222_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8397__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8810_ _1497_ _3181_ _3963_ _3939_ _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9133__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8741_ _3908_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4958__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5953_ _1309_ _1340_ _1342_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6524__B _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5080__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _0319_ _0332_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5884_ as2650.stack\[3\]\[0\] _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8672_ as2650.stack\[6\]\[3\] _3860_ _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _2875_ _2876_ _2675_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4835_ _4314_ _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6175__A4 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7554_ net34 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5383__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _4359_ _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _1818_ _1819_ _1821_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7485_ _2711_ _2696_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4697_ _4262_ _4289_ _4290_ _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8321__A2 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5135__A2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6332__A1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6436_ _0413_ _1751_ _1758_ _0666_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9155_ _0252_ clknet_leaf_71_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6367_ _4372_ _1467_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_103_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8106_ _3278_ _3336_ _3327_ _3282_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5318_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9086_ _0183_ clknet_leaf_23_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6298_ _1634_ _1635_ _1636_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8037_ _2527_ _3269_ _1687_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5249_ _4165_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8388__A2 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6399__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7060__A2 _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8939_ _0050_ clknet_leaf_58_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4949__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7899__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8808__C _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4908__I _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6626__A2 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4637__A1 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8824__B _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7051__A2 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5062__A1 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4643__I _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8000__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8551__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _4144_ _4213_ _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6562__A1 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5365__A2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4551_ as2650.r123\[1\]\[1\] as2650.r123\[0\]\[1\] as2650.r123_2\[1\]\[1\] as2650.r123_2\[0\]\[1\]
+ _4066_ _4062_ _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5474__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8303__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7270_ _2529_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4482_ _4075_ _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6314__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5117__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6221_ _1554_ _1566_ _1567_ _1568_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6865__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8785__I _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4876__A1 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8067__A1 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6152_ _0468_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8067__B2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _0513_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7814__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7814__B2 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ as2650.stack\[0\]\[6\] _1445_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5034_ _4320_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5649__I as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6985_ _2289_ _2282_ _2290_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4553__I _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8790__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8724_ _3898_ _3899_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4800__A1 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8655_ as2650.stack\[7\]\[11\] _3851_ _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5867_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8542__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7606_ _2848_ _2852_ _2859_ _2607_ _1588_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4818_ _4271_ as2650.cycle\[10\] _4412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5356__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8586_ as2650.psu\[5\] _3700_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7537_ _2773_ _2738_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4749_ _4244_ _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6305__A1 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7468_ net55 _2601_ _2723_ _2724_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net51 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7813__B _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput25 net25 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6419_ _0397_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput36 net36 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7399_ _4336_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8058__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9138_ _0235_ clknet_leaf_44_wb_clk_i as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7805__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6608__A2 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9069_ _0166_ clknet_leaf_50_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7104__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__A1 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8230__A1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7033__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5044__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8781__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6792__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6139__A4 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8297__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__A1 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8049__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__C _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8049__B2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__I _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7272__A2 _4439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7949__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4625__A4 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8221__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5469__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5035__B2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6770_ _2084_ _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7980__B1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5721_ as2650.stack\[7\]\[14\] _1043_ _1044_ as2650.stack\[6\]\[14\] _1047_ _1125_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8524__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8440_ _1416_ _3633_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5652_ _0917_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _4134_ _4196_ _4167_ _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8371_ _3000_ _3563_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5583_ _0988_ _0540_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7322_ _2524_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8288__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4534_ _4127_ _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7253_ _4283_ _4348_ _0556_ _1520_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4465_ _4058_ _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5932__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8448__C _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6302__A4 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6204_ _1529_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7184_ _0706_ as2650.psu\[1\] _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4548__I _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6135_ _1095_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7263__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8460__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _1436_ _1347_ _1352_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A1 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _0429_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8183__C _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8212__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__C _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A1 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6968_ as2650.r123_2\[2\]\[7\] _1856_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8707_ _0468_ _3884_ _3886_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ _1312_ _1273_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6899_ _0740_ _1812_ _2198_ _2211_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7527__C _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8638_ as2650.stack\[7\]\[5\] _3841_ _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8569_ _1303_ _3727_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8279__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__C _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6829__A2 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5888__I0 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__A2 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8451__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5568__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8506__A2 _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4921__I as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7437__C _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7565__I0 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__I1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7245__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8442__A1 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8442__B2 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7679__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _3170_ _1678_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7871_ _2673_ _1525_ _3117_ _1252_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5199__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8745__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6822_ _2122_ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6756__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5559__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _2019_ _2031_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4831__I _4424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ as2650.stack\[1\]\[13\] _0704_ _0710_ as2650.stack\[0\]\[13\] _1109_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6684_ _1964_ _1994_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8423_ _3433_ _1049_ _3344_ _3627_ _2781_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7181__A1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8354_ _2816_ _3577_ _3313_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _0905_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5731__A2 _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8459__B _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7305_ _0660_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4479__S _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4517_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _4110_ _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8285_ _3194_ _3502_ _3510_ _0435_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5497_ as2650.psu\[2\] _0713_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7236_ _0317_ _4340_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8681__A1 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7167_ as2650.r123_2\[0\]\[4\] _2437_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7236__A2 _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8433__A1 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _0737_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7098_ _1216_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ as2650.pc\[13\] _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6995__A1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8736__A2 _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5837__I _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__I _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7172__A1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5722__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8121__B1 _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7475__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6278__A3 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8424__A1 _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5238__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8727__A2 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7448__B _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__A4 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5410__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8123__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6578__I _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _0594_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8663__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8070_ _3246_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5282_ _0544_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ as2650.r123_2\[1\]\[4\] _2306_ _2317_ _2310_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__A2 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8415__A1 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5229__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8972_ _0083_ clknet_leaf_15_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8718__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7854_ _2511_ _2517_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6805_ _2078_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7785_ _3026_ _3034_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4997_ _0419_ _0325_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6736_ _0791_ _2048_ _1818_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ _4160_ _1859_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7154__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8351__B1 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7154__B2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8406_ _3626_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _0683_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5704__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6901__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6598_ _1882_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8337_ _1390_ _3560_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5549_ _0951_ _0522_ _0955_ _0668_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7457__A2 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0__f_wb_clk_i clknet_0_wb_clk_i clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8654__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8268_ _3263_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7219_ _0465_ _4051_ _2480_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_132_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8199_ as2650.stack\[3\]\[5\] _3246_ _1573_ as2650.stack\[2\]\[5\] _3427_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4691__A2 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8709__A2 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7393__A1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7782__I _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8893__A1 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7731__B _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__B1 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7620__A2 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7957__I _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ _4354_ _4246_ _0345_ _0294_ _0346_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ _4432_ _4365_ _4437_ _4443_ _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7384__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8581__B1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ _2544_ _2820_ _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4782_ _4375_ _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _0676_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7136__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9240_ net48 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6452_ _1420_ _1772_ _1778_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5698__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9062__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _4358_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9171_ _0268_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6383_ _1654_ _1720_ _1704_ _1467_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5162__A3 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8122_ _3316_ _3318_ _3342_ _3352_ _3220_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7439__A2 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8053_ _3283_ _3284_ _4448_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ net7 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6111__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5940__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _2038_ _1924_ _2304_ as2650.r123_2\[1\]\[0\] _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5196_ _0584_ _0595_ _0600_ _0603_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_84_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8955_ _0066_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7906_ _0313_ _0327_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8886_ _3185_ _4030_ _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4976__A3 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7837_ _3083_ _3084_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7375__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6178__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7768_ _2940_ _2966_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6719_ _1998_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7699_ _2882_ _2938_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8324__B1 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8875__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7107__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__A3 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8627__A1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7850__A2 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4664__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5861__A1 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4466__I _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7602__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7777__I _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__A1 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6169__A2 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8563__B1 _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7669__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8866__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8866__B2 _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8922__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _0433_ _0458_ _0459_ _0467_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5852__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5604__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8740_ _3907_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ as2650.stack\[2\]\[4\] _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5080__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4903_ _0321_ _4350_ _0328_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_52_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8671_ _2287_ _3859_ _3863_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7357__A1 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5883_ _1271_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7622_ _1322_ _2583_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4834_ _4258_ _4427_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7553_ _2346_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _4358_ _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6580__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6504_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8857__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7484_ net33 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ as2650.halted _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _1767_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5135__A3 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6332__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9154_ _0251_ clknet_leaf_44_wb_clk_i as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6366_ _4387_ _0620_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4894__A2 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8105_ _2664_ _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ as2650.stack\[1\]\[8\] _0725_ _0726_ as2650.stack\[0\]\[8\] _0727_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_9085_ _0182_ clknet_leaf_23_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _1473_ _0483_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8036_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7832__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _0655_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4646__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7596__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__A2 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8938_ _0049_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8869_ _1192_ _1193_ _1208_ _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7899__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__B _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8848__A1 _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7520__A1 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8945__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6323__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5677__A4 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__A2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7823__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5513__C _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4637__A2 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A1 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4924__I _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5062__A2 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6344__C _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8000__A2 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6011__A1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6562__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4550_ _4143_ _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ as2650.r0\[7\] _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6314__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6220_ _1507_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4876__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _1487_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_41_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ as2650.r123\[3\]\[7\] _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9100__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _1317_ _1444_ _1447_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5033_ _0451_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ as2650.stack\[5\]\[3\] _2283_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7210__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8723_ _3892_ _2317_ _3893_ _1039_ _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5935_ _1211_ _1306_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8527__B1 _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4800__A2 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8654_ _1792_ _3848_ _3853_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5866_ _4343_ _1257_ _1263_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7605_ _2854_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4817_ as2650.addr_buff\[7\] _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8585_ _0355_ _1078_ _3796_ _3797_ _3693_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8968__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _1191_ _1184_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8041__I _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7536_ _2766_ _1021_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4564__A1 _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _4341_ _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7467_ _4431_ _1710_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ _4263_ _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7502__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6305__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6418_ _0736_ _1215_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput15 net15 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput26 net26 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ _2647_ _2655_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput37 net37 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9137_ _0234_ clknet_leaf_53_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6349_ _1660_ _1648_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7805__A2 _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6608__A3 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9068_ _0165_ clknet_leaf_59_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5816__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8019_ _3241_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7569__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6792__A2 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__B2 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8297__A2 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9123__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__A2 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__I as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8049__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5283__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__I _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8221__A2 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7980__A1 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7980__B2 _4327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ as2650.stack\[5\]\[14\] _0705_ _0711_ as2650.stack\[4\]\[14\] _1124_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5651_ as2650.holding_reg\[5\] _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ _4192_ _4195_ _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8370_ _3188_ _3592_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5582_ _4118_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7321_ _2526_ _2579_ _2580_ _1568_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ as2650.r0\[3\] _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8288__A2 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__A1 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7252_ _0310_ _2494_ _1749_ _4290_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_105_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ as2650.ins_reg\[0\] _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6203_ _1530_ _1552_ _1553_ _1549_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4829__I _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7183_ _2453_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6134_ _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7799__B2 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7263__A3 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8460__A2 _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _0707_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5016_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8748__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8036__I _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8212__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6223__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _2038_ _2276_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7971__A1 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8706_ _0480_ _0570_ _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5918_ _1314_ _1306_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6898_ as2650.r123_2\[2\]\[4\] _1856_ _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8637_ _2291_ _3840_ _3842_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5849_ _0396_ _1248_ _1249_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__9146__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _3731_ _3781_ _3782_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7519_ _2701_ _2774_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8279__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8499_ _4400_ _4318_ _3343_ _1638_ _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_107_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5888__I1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8203__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6214__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__B _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7025__I _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4551__I1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7245__A3 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__A2 _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9240__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8284__C _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9019__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ _0386_ _0442_ _0361_ _0454_ _0303_ net27 _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6821_ _2124_ _2135_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6756__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _2066_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5703_ _0748_ _1078_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _1999_ _1993_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7705__A1 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6508__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8422_ _3632_ _3640_ _4368_ _3642_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5634_ as2650.stack\[3\]\[12\] _0714_ _0710_ as2650.stack\[0\]\[12\] _1040_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8353_ _3433_ _0832_ _3426_ _3562_ _3576_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_129_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5565_ as2650.stack\[1\]\[11\] _0725_ _0726_ as2650.stack\[0\]\[11\] _0718_ as2650.stack\[2\]\[11\]
+ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_129_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7304_ _2560_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4516_ _4109_ _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8284_ _1328_ _4415_ _3509_ _0813_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__8130__A1 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5496_ as2650.stack\[3\]\[10\] _0821_ _0822_ as2650.stack\[2\]\[10\] _0904_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7235_ _2492_ _2494_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4559__I _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5495__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8418__C1 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7166_ _2209_ _2406_ _2416_ _2439_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4495__S _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _0572_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8433__A2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _1659_ _2363_ _2383_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6048_ _1387_ _1420_ _1421_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7999_ _3132_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7944__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__I _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5707__B1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5183__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8121__A1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8121__B2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4469__I _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6278__A4 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8188__A1 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7935__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4932__I _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8360__A1 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _0607_ _0619_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8112__A1 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8663__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5281_ _0661_ _0665_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7020_ _1921_ _1934_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7871__B1 _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7911__C _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6426__B2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8971_ _0082_ clknet_leaf_15_wb_clk_i net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7922_ _1802_ _3162_ _0530_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5003__I _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8179__A1 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7853_ _4222_ _1482_ _0557_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4842__I _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6804_ _2088_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7784_ _1400_ _2728_ _3031_ _3033_ _0305_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4996_ _0323_ _0403_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _4218_ _1837_ _2050_ _2047_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _1942_ _1981_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8351__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8351__B2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8405_ _1416_ _3625_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5617_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5165__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ _4139_ _1895_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8336_ _1379_ _3530_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5548_ _4212_ _0554_ _0954_ _0521_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8103__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_opt_3_0_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_opt_3_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8267_ _3378_ _3462_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8654__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _4156_ _0879_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6665__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7218_ _2478_ _2479_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8198_ _3343_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7149_ _2061_ _2419_ _2420_ _2425_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6968__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6009__I _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4752__I _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8590__A1 _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7393__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout50 net51 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8342__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8893__A2 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4903__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__A1 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__A2 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6408__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6408__B2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__A3 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7459__B _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7908__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4662__I _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4850_ _4440_ _4442_ _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7384__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8581__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8581__B2 _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A1 as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ as2650.ins_reg\[3\] as2650.ins_reg\[2\] _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7973__I _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6520_ _1813_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8333__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7136__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ as2650.stack\[0\]\[12\] _1774_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__A1 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6344__B1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _0748_ _0775_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_127_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9170_ _0267_ clknet_leaf_5_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5426__C _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6382_ _1711_ _1715_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8121_ _3344_ _3327_ _3351_ _3258_ _2816_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _0742_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7439__A3 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8636__A2 _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6647__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ _0784_ _4151_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7641__C _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5264_ _4209_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__B _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7003_ _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4837__I _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5195_ _4193_ _4376_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_68_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7072__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8954_ _0065_ clknet_leaf_33_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7905_ _3138_ _3149_ _3150_ _2629_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8885_ _3184_ _4028_ _1212_ _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4976__A4 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7836_ as2650.pc\[12\] _1142_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7375__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7767_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4979_ _4273_ as2650.cycle\[1\] _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6583__B1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6718_ _2002_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7698_ _2857_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8324__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8324__B2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__A1 _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ _1946_ _1957_ _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8875__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6886__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8319_ _2329_ _4436_ _3543_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5352__B _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__I _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4664__A3 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7063__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7994__S _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4482__I _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8563__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8563__B2 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7118__A2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__A1 as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6877__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4657__I _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _1333_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ as2650.cycle\[1\] _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8670_ as2650.stack\[6\]\[2\] _3860_ _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5882_ _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8554__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7621_ _2860_ _2874_ _2673_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4833_ _4355_ _4408_ _4422_ _4426_ _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_33_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7552_ _2796_ _2801_ _2802_ _2806_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4764_ _4357_ _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7109__A2 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _0367_ _0301_ _1816_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7483_ _2735_ _2738_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4695_ _4267_ _4275_ _4286_ _4288_ _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7208__I _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _1674_ _1751_ _1758_ _0494_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6332__A3 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9153_ _0250_ clknet_leaf_45_wb_clk_i as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5540__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _0882_ _4192_ _1089_ _1143_ _4215_ _0675_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__8609__A2 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5951__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5540__B2 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8104_ _1287_ _3279_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ _0709_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9084_ _0181_ clknet_leaf_23_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7371__C _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _4319_ _1459_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8035_ _3216_ _3218_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8039__I _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _0656_ _0533_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5178_ _4160_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A1 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6782__I _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__A1 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8937_ _0048_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__I _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8868_ _0485_ _1631_ _3990_ _4016_ _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__8545__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8545__B2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7819_ _2526_ _3066_ _3067_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7899__A3 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8799_ _3952_ _0502_ _1248_ _1476_ _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7520__A2 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5531__B2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__A1 _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7788__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__B _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8784__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7339__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8536__A1 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7737__B _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__I _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5770__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A2 _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5770__B2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4480_ _4072_ _4073_ _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _1477_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7275__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _0512_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ as2650.stack\[0\]\[5\] _1445_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5032_ _0353_ _4349_ _0320_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_81_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_81_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7027__A1 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _1299_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8722_ as2650.r123\[1\]\[4\] _3890_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _1328_ _1306_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8527__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8527__B2 _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8653_ as2650.stack\[7\]\[10\] _3851_ _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5865_ _4246_ _1265_ _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_80_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7604_ _2855_ _2857_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4816_ _4409_ _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__C _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _1189_ _1190_ _1185_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8584_ _3688_ _1086_ _0354_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7535_ _1313_ _1091_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4747_ _4226_ _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4564__A2 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7466_ _4435_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4678_ _4271_ as2650.cycle\[12\] _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6417_ _1750_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5513__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5681__I _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _2639_ _2561_ _2652_ _2654_ _2612_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xoutput16 net16 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput38 net38 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9136_ _0233_ clknet_leaf_53_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6348_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9067_ _0164_ clknet_leaf_52_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8463__B1 _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6608__A4 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6279_ _1616_ _1617_ _1210_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8018_ _1572_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7569__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8766__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6241__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4760__I _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8912__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5077__B _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8049__A3 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8835__C _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4935__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7311__I _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8221__A3 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7980__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9238__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5650_ _4116_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _4155_ _4194_ _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5581_ _0984_ _0985_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5743__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _2541_ _2525_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4532_ _4125_ _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7914__C _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7496__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7251_ _1643_ _1266_ _2509_ _0475_ _2510_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6299__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6543__I0 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4463_ _4056_ _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ net45 _1538_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ as2650.r123_2\[0\]\[7\] _2437_ _2452_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7248__A1 _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9098__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _1478_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _1387_ _1434_ _1435_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7263__A4 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8460__A3 _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4845__I _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6471__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8212__A3 _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8935__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6966_ _2250_ _2260_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7971__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8705_ _3884_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6897_ _1830_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8636_ as2650.stack\[7\]\[4\] _3841_ _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _4358_ _0390_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8567_ _0969_ _3750_ _3038_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5779_ as2650.r123\[0\]\[7\] _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7518_ _2633_ _2659_ _2702_ _2704_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8498_ _2821_ _3712_ _3713_ _3715_ _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7487__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7449_ _2703_ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6534__I0 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6300__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7239__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9119_ _0216_ clknet_leaf_80_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8227__I _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__I _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__I _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8739__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A1 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7411__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6970__I _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__I as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7478__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7306__I _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6150__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8846__B _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4551__I2 as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4665__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__A2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__I _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _2021_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6751_ _1120_ _2005_ _2016_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ _0644_ _1086_ _1106_ _0913_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6682_ _1966_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7705__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8421_ _2473_ _3636_ _3641_ _3455_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5633_ _0748_ _1009_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8352_ _3571_ _3574_ _3575_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5564_ _0970_ _0818_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7469__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7303_ _1752_ _0660_ _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4515_ _4108_ _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8283_ _2585_ _2884_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5495_ as2650.stack\[5\]\[10\] _0725_ _0726_ as2650.stack\[4\]\[10\] _0825_ _0903_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7216__I _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8130__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7234_ _4387_ _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6141__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7660__B _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6692__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7165_ _2421_ _2414_ _2411_ _1303_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _0446_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7096_ _2382_ _2359_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7641__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6047_ as2650.stack\[1\]\[12\] _1397_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7886__I _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9113__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7998_ _2362_ _3140_ _3229_ _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4758__A2 _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5955__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _2251_ _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8619_ _2385_ _0678_ _1615_ _1139_ _3730_ _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_127_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8121__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A1 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7570__B _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7880__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A1 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5802__C _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4485__I _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7796__I _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8188__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7935__A2 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5946__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6205__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A1 _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__I _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _0669_ _0673_ _0687_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8576__B _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8663__A3 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7871__A1 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7871__B2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8970_ _0081_ clknet_leaf_15_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5634__B1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7921_ _1463_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _2526_ _3098_ _3099_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6803_ _1954_ _2021_ _2072_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5937__A1 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7783_ _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4995_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _0786_ _2049_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ as2650.r0\[7\] _1869_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8330__I _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8404_ _1406_ _3602_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5616_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5165__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _1910_ _1911_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8335_ _3558_ _3559_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _0953_ _0554_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6114__A1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8266_ _3488_ _3489_ _3492_ _1047_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5478_ _0880_ _0522_ _0885_ _0668_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6785__I _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7217_ _0341_ _1468_ _0481_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8197_ _3424_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A1 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7148_ _2421_ _2422_ _2423_ _1540_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_86_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7079_ as2650.addr_buff\[2\] _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4979__A2 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout51 net14 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8342__A2 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5085__B _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__A2 _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6105__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8396__B _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__A1 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6408__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5104__I as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7081__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4943__I _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8030__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5919__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8581__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4780_ _4373_ _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_35_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8333__A2 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8150__I _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _1414_ _1771_ _1777_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5147__A2 _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5401_ _0580_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6381_ as2650.overflow _1718_ _1500_ as2650.psl\[5\] _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8097__A1 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5332_ _0575_ _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8120_ _3350_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7844__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8051_ net7 _4161_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6647__A2 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5263_ _0609_ _0672_ _0612_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__C _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7002_ _1633_ _1829_ _1854_ _0322_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5194_ as2650.holding_reg\[0\] _0591_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5014__I _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7072__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8953_ _0064_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7904_ net52 _3138_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8884_ _4029_ _4031_ _3647_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7835_ _3018_ _3080_ _3082_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8572__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7766_ as2650.pc\[9\] _1378_ _2840_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5386__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ _0387_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6583__B2 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6717_ _2007_ _2033_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _2853_ _2881_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8324__A2 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__I _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6648_ _1947_ _1956_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5138__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6886__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8318_ _2361_ _2891_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8249_ _1321_ _0410_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4664__A4 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7063__A2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8235__I _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__I _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8563__A2 _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6574__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A2 as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__A1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8079__A1 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A1 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8251__A1 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5950_ _1333_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8003__A1 _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5881_ _0698_ _1273_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8554__A2 _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7620_ _4362_ _2861_ _2872_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_33_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _4363_ _4366_ _4425_ _4426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7551_ _2685_ _2805_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4763_ _4356_ _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _0566_ _1808_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7482_ _2701_ _2705_ _2737_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4694_ _4232_ _4250_ _4287_ _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _0615_ _1761_ _1759_ _1766_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4879__A1 _4433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9152_ _0249_ clknet_leaf_46_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6364_ _4414_ _0672_ _1561_ _1094_ _4189_ _1022_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5540__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7817__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8103_ _0436_ _3333_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5315_ _0703_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9083_ _0180_ clknet_leaf_22_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6295_ _1633_ _1622_ _1469_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8034_ _3220_ _3266_ _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8490__A1 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5246_ _0532_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5177_ _0539_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A2 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8936_ _0047_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8867_ _1626_ _4015_ _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7818_ _3049_ _2786_ _3038_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8798_ _4248_ _0368_ _1264_ _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7749_ as2650.pc\[10\] _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8481__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6973__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8233__A1 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8784__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8991__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8536__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4558__B1 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8839__A3 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A3 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__I _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ as2650.r123\[3\]\[6\] _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7275__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _1309_ _1444_ _1446_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8472__A1 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _0383_ _4370_ _0303_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__A1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7027__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _2287_ _2282_ _2288_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6786__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8721_ _0967_ _3883_ _3897_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5933_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8527__A2 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8652_ _1789_ _3848_ _3852_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6538__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ _4358_ _0556_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _1313_ _1500_ _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4815_ _4333_ _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8583_ _3734_ _1104_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5795_ _1195_ _1196_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5210__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6123__I _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7534_ _2788_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ _4336_ _4339_ _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4564__A3 as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7465_ _2721_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4677_ _4264_ _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5962__I _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6416_ _0342_ _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6710__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _2561_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6279__B _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput17 net17 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9135_ _0232_ clknet_leaf_56_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6347_ _0350_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8463__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9066_ _0163_ clknet_leaf_51_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _1120_ _1087_ _1017_ _0949_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__8463__B2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5277__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8017_ _2387_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5229_ _0330_ _0325_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8215__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6777__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5202__I _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7838__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8919_ _0030_ clknet_leaf_35_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8518__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8513__I _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6529__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7129__I _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8151__B1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4488__I _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5268__A1 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6409__S _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8757__A2 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5112__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4951__I _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _4171_ _4193_ _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5580_ _0984_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4531_ _4124_ _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7250_ _0483_ _1278_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6299__A3 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ _4053_ _4055_ _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6543__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6201_ _0969_ _1533_ _1551_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7181_ _2272_ _2406_ _2415_ _2451_ _2416_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7248__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _1462_ _1464_ _1486_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8445__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ as2650.stack\[1\]\[14\] _1369_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _4288_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8748__A2 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6118__I _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5022__I _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__B _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _2273_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5431__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8704_ _0741_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ as2650.pc\[5\] _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _2199_ _2208_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8635_ _3833_ _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _0494_ _0630_ _4316_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8566_ _3769_ _3779_ _3780_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5778_ _1119_ _0983_ _1181_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6931__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7517_ _2766_ net11 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4729_ _4322_ _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8497_ _1764_ _3714_ _2341_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7448_ _2634_ _2636_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7487__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ _2634_ _2636_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7239__A2 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8436__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9118_ _0215_ clknet_leaf_80_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9049_ _0004_ clknet_leaf_29_wb_clk_i as2650.cycle\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9192__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8739__A2 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__I _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7411__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7568__B _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5867__I _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4771__I _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7287__C _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7175__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5725__A2 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__C _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8427__A1 _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4551__I3 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7322__I _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6989__A1 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _0777_ _2003_ _2014_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ _1016_ _1101_ _1105_ _0644_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6681_ _1961_ _1996_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7166__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8420_ _3175_ _3627_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ _0644_ _1015_ _1037_ _0913_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7961__I0 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8351_ _2728_ _3566_ _3562_ _0557_ _4443_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__9065__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5563_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8115__B1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7302_ _2561_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7469__A2 _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ _4061_ _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8666__A1 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8282_ _3503_ _3504_ _3507_ _0723_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_5494_ as2650.stack\[7\]\[10\] _0821_ _0822_ as2650.stack\[6\]\[10\] _0902_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7233_ _0550_ _0561_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6141__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5017__I _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8418__A1 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8418__B2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7164_ _1049_ _2428_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ _1466_ _1469_ _0736_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7095_ _0532_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7641__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6292__B _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5687__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7997_ _3222_ _2596_ _0463_ _2329_ _0814_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _2254_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_41_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _1017_ _2156_ _2167_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8618_ _3827_ _3828_ _1699_ _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6365__C1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5707__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6904__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8549_ _3202_ _3764_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8106__B1 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6311__I _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7851__B _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A2 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7880__A2 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4694__A2 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4766__I _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__I _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__C _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5643__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__B _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8593__B1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5946__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9088__CLK clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7148__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8345__B1 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7148__B2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8925__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7320__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4685__A2 _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8148__I _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8820__A1 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7987__I _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7920_ _0490_ _0497_ _0369_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7851_ net53 _2786_ _3038_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _1186_ _2005_ _2073_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_64_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7782_ _2336_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4994_ _4409_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5937__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6733_ _1813_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7139__A1 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6664_ _4098_ _1872_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8403_ _3069_ _3499_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5615_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6595_ _1905_ _1910_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8334_ _1381_ _3269_ _3354_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8639__A1 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5546_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8265_ as2650.stack\[7\]\[6\] _3250_ _3251_ as2650.stack\[6\]\[6\] _3491_ _3492_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_117_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _0883_ _0682_ _0884_ _0685_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8486__C _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7216_ _1246_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8196_ _2789_ _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A2 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7147_ _0832_ _2409_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7614__A2 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8811__A1 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7078_ _1718_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_5__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8811__B2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5625__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ as2650.stack\[1\]\[10\] _1397_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_5_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7846__B _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout52 net26 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A2 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8521__I _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8878__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8948__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7550__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6105__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__A2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A1 _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4496__I _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8802__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7369__A1 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8030__A2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_90 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_127_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7541__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _0797_ _0803_ _0807_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6380_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_75_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_75_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8587__B _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5331_ _0551_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8097__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9103__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8050_ _3281_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7844__A2 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__C _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5262_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _0601_ _0599_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__A1 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8952_ _0063_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7903_ _3144_ _3147_ _3148_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8883_ _3191_ _4030_ _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6126__I _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7834_ _3041_ _3016_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7765_ _3014_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4977_ _4444_ _0389_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5965__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7780__A1 _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__A2 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6716_ _2010_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4594__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7696_ _0441_ _2947_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ _0988_ _1906_ _1944_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6578_ _1871_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8497__B _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8317_ _2362_ _3541_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8088__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _0616_ _0853_ _0925_ _0926_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _0397_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8179_ _3402_ _3407_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5205__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6271__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8548__B1 _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5875__I _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7771__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9126__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8787__B1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8426__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8251__A2 _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ as2650.cycle\[2\] _4265_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8003__A2 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5880_ _1277_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _4424_ _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7762__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8161__I _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7550_ _1094_ _1086_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4576__A1 as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ as2650.cycle\[6\] _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6501_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7481_ _2710_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7514__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _4277_ _4240_ _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6432_ _0348_ _1764_ _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__A2 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9151_ _0248_ clknet_leaf_53_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6363_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8102_ _4050_ _3332_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5314_ as2650.stack\[6\]\[8\] _0719_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9082_ _0179_ clknet_leaf_22_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7817__A2 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ _1632_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5828__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ _2527_ _3221_ _3265_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5245_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8490__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5176_ _0584_ _4164_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4864__I _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8242__A2 _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7045__A3 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6253__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8935_ _0046_ clknet_leaf_57_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8866_ _0489_ _3951_ _3940_ _4402_ _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6005__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7817_ _1409_ _2530_ _3065_ _2996_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8797_ _3168_ _0739_ _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7753__A1 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8071__I _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7748_ _2787_ _2997_ _2998_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7679_ net37 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7505__A1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6308__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7415__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5819__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6492__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7744__A1 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7744__B2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4558__A1 _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8839__A4 _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7753__C _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7325__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8472__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5030_ _4437_ _0381_ _0446_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8224__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6981_ as2650.stack\[5\]\[2\] _2283_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7983__A1 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ as2650.pc\[7\] _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8720_ _3885_ _2314_ _3888_ as2650.r123\[1\]\[3\] _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8651_ as2650.stack\[7\]\[9\] _3851_ _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5863_ _1131_ _0367_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7735__A1 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7602_ _2766_ net11 _1091_ _2788_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__A1 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _4363_ _4366_ _4407_ _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8582_ _1508_ _3783_ _3795_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5794_ _1195_ _1196_ _0616_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5210__A2 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7533_ as2650.pc\[5\] _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4745_ _4338_ _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7464_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4676_ _4269_ _4255_ _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6415_ _1676_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7395_ _2650_ _2651_ _2649_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6710__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9134_ _0231_ clknet_leaf_56_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput29 net29 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6346_ _1589_ _1613_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9065_ _0162_ clknet_leaf_49_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _0876_ _0777_ _0662_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8463__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8016_ as2650.stack\[1\]\[0\] _3242_ _3245_ as2650.stack\[0\]\[0\] _3248_ _3249_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5228_ _0583_ _0635_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_131_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5159_ _0545_ _0548_ _0554_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__9102__D _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5029__A2 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6777__A2 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A1 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8918_ _0029_ clknet_3_1__leaf_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__A1 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8849_ _3996_ _3999_ _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6529__A2 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__B2 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5201__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4960__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__I _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5268__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4718__B _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8206__A2 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__A1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8704__I _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4779__A1 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5440__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__B _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8390__A1 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8579__C _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4530_ _4119_ _4121_ _4123_ _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__8142__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4461_ _4054_ _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8693__A2 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6200_ _1550_ _1535_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7180_ _1211_ _2409_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _1471_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8445__A2 _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5013_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6964_ _2254_ _2258_ _2255_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5431__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8703_ _1633_ _1132_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5459__B _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1088_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7708__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6895_ _2057_ _2206_ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7708__B2 _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6134__I _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8634_ _3833_ _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5846_ as2650.halted _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7184__A2 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5195__A1 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _1123_ _1130_ _0745_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8565_ _2373_ _3754_ _0426_ _1550_ _4212_ _2606_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__6931__A2 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__C _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7516_ _2722_ _2742_ _2771_ _0441_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4728_ _4238_ _4169_ _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8496_ _4057_ _0493_ _4359_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7447_ _1292_ _1717_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7487__A3 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8684__A2 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4659_ _4252_ _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7378_ _2635_ _2623_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9117_ _0214_ clknet_leaf_80_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6329_ _4185_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8436__A2 _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__A1 as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9048_ _0003_ clknet_leaf_14_wb_clk_i as2650.cycle\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7568__C _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8372__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7175__A2 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8372__B2 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5883__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8399__C _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8124__A1 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__I _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6438__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_29_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4962__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ _1016_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _1963_ _1995_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8363__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _1016_ _1031_ _1036_ _0808_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7961__I1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8350_ _3281_ _3562_ _3573_ _3234_ _2548_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5562_ _0949_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8115__B2 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7301_ _2560_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4513_ _4106_ _4078_ _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8281_ as2650.stack\[7\]\[7\] _2389_ _3380_ as2650.stack\[4\]\[7\] _3506_ _3507_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_5493_ _0866_ _0900_ _0580_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7232_ _4348_ _4284_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7163_ _2404_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8418__A2 _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6429__A1 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ _1467_ _1468_ _0495_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7094_ _1502_ _2363_ _2381_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ as2650.r123\[0\]\[4\] _1374_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7669__B _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7929__A1 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5968__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4872__I _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7996_ _2715_ _2539_ _3228_ _0399_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6947_ _2255_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8354__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _2164_ _2166_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8617_ _2230_ _0503_ _3508_ _0733_ _3770_ _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6365__B1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5829_ _0671_ _1010_ _1226_ _0892_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6365__C2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8548_ _1545_ _3750_ _3753_ _3763_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8106__A1 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8106__B2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8657__A2 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8479_ _1632_ _0368_ _1264_ _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6668__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__A3 _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5891__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7093__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6039__I _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8290__B1 _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6840__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4782__I _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8593__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8593__B2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8345__A1 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8345__B2 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5159__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8648__A2 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5331__A1 _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7333__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8281__B1 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7850_ _3069_ _2530_ _3097_ _2996_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8584__A1 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _2068_ _2091_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7781_ _3000_ _2597_ _2331_ _3030_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4993_ _0384_ _0402_ _0409_ _0416_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6732_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6663_ _1977_ _1978_ _1979_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8402_ _3621_ _3623_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5614_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9182__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6594_ _0776_ _1902_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5545_ net10 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8333_ _3316_ _3532_ _3550_ _3557_ _3220_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5028__I _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8264_ _3490_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5476_ _4214_ _0683_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6114__A3 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7215_ _2475_ _2476_ _2477_ _1568_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4867__I _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8195_ _1304_ _1296_ _3356_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7146_ _2411_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7077_ _2365_ _2360_ _2368_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8811__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5625__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8575__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8007__C _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7979_ _3211_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8327__B2 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout53 net41 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8878__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7550__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4777__I _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7853__A3 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5864__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8263__B1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6813__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9055__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_80 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_91 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_127_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8318__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7328__I _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _0737_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7000_ _1633_ _1829_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5192_ _0591_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7057__A1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8951_ _0062_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7902_ _0309_ _1749_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8882_ _1732_ _3190_ _4028_ _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7833_ _1406_ _1142_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7764_ _1399_ _1141_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8309__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4976_ _0394_ _4366_ _0395_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7780__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ _2017_ _2019_ _2031_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_7695_ _2666_ _2933_ _2945_ _2946_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7238__I _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6142__I _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6646_ _1938_ _1959_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5138__A4 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6577_ _1879_ _1884_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8316_ _2891_ _3540_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5528_ _0925_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7296__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__I _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8247_ _1321_ _3442_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _4148_ _4154_ _4164_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9105__D _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8178_ _3128_ _3403_ _3406_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9078__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7048__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ _0737_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6317__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8548__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8915__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4585__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6987__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8200__C _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7287__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8787__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8787__B2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6227__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_2_0_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__I _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7211__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _4423_ _4424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7762__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _4331_ _4352_ _4354_ _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4576__A2 as2650.alu_op\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5773__B2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _0630_ _4307_ _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7480_ net10 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4692_ _4276_ _4280_ _4281_ _4285_ _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7514__A2 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5525__A1 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6431_ _0348_ _1502_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6722__B1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9150_ _0247_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6362_ _4306_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8110__C _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8101_ _4429_ _3324_ _3331_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5313_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9081_ _0178_ clknet_leaf_22_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6293_ _1465_ _0476_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ _0532_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8032_ _3233_ _3240_ _3256_ _3258_ _3264_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4500__A2 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5175_ _4394_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8778__A1 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7450__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6253__A2 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8934_ _0045_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5041__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8865_ _4008_ _4013_ _4014_ _0349_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_73_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7816_ _2814_ _3054_ _3064_ _2961_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8796_ _3947_ _3949_ _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4813__C _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7747_ _2978_ _2829_ _2830_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ as2650.cycle\[4\] _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7678_ _2686_ _2923_ _2928_ _2929_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8702__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5516__A1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ _1944_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7269__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6492__A2 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5886__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8865__C _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7341__I _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8881__B _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _1293_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5931_ _1302_ _1325_ _1326_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8650_ _3846_ _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _0474_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7735__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7601_ _2792_ _2790_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4549__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ _4368_ _4326_ _4404_ _4406_ _4407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8581_ _2144_ _0426_ _1589_ _3786_ _3794_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5793_ _1173_ _1170_ _1163_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _2786_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4744_ as2650.cycle\[2\] _4337_ _4271_ _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7499__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7463_ _4434_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4675_ _4268_ _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_107_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6414_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6171__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7394_ _2649_ _2650_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 net19 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_127_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9133_ _0230_ clknet_leaf_46_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7960__B _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6345_ _1615_ _1621_ _1648_ _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4721__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9064_ _0161_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6276_ _1489_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7671__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4875__I _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6474__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5227_ _0636_ _0605_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8015_ _3247_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5158_ _0555_ _0559_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8791__B _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7423__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6226__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8620__B1 _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _0506_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9116__CLK clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8917_ _0028_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5985__A1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8848_ _3997_ _3998_ _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8779_ as2650.stack\[4\]\[7\] _3932_ _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8151__A2 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6162__A1 _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4785__I _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7662__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4476__A1 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7414__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7414__B2 _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__A2 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7717__A2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8142__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4460_ as2650.alu_op\[1\] _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _1475_ _1476_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7653__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ as2650.r123\[0\]\[6\] _1374_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9139__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5012_ _4290_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _2251_ _2259_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8702_ _1800_ _3874_ _3882_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6415__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5914_ _1302_ _1309_ _1311_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6894_ _1015_ _1826_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7708__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5719__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8633_ _2289_ _3834_ _3839_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5845_ _1246_ _0347_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_107_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8381__A2 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5195__A2 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8564_ _3755_ _3776_ _3778_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5776_ _1133_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7515_ _2600_ _2769_ _2770_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4727_ _4311_ _4314_ _4320_ _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8495_ _1493_ _4314_ _1531_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7446_ _2701_ _2702_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4658_ as2650.ins_reg\[3\] _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8684__A3 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7892__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7377_ as2650.pc\[1\] _0784_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _4104_ _4168_ _4182_ _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9116_ _0213_ clknet_3_6__leaf_wb_clk_i as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _1561_ _1099_ _4199_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7644__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9047_ _0002_ clknet_3_2__leaf_wb_clk_i as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6259_ _0848_ _0853_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8805__I _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5958__A1 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8124__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4697__A1 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7635__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8832__B1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__I _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5949__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6235__I _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_69_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_69_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7775__B _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8363__A2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _1016_ _1035_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8115__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7300_ _4430_ _1531_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ _4105_ _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5492_ _0890_ _0896_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8280_ _3505_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7231_ _2484_ _2490_ _2491_ _1689_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7874__A1 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ _2436_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _4316_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6429__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7093_ _2380_ _2367_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _1416_ _1391_ _1372_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8625__I _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7929__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ _1276_ _0392_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6145__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _2182_ _2183_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _2180_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8616_ as2650.psu\[7\] _3772_ _1460_ _3826_ _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6365__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _0941_ _1224_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6365__B2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8547_ _4214_ _0466_ _3730_ _3762_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4915__A2 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5759_ _1161_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__S0 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8478_ _1541_ _3695_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7865__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6668__A2 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7429_ _4339_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5340__A2 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7617__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8290__A1 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7093__A2 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8290__B2 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A1 _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8042__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7856__A1 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7608__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8281__B2 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6393__C _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8033__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8971__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6800_ _2071_ _2090_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7780_ _3027_ _3011_ _3028_ _3029_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4992_ _0413_ _4366_ _0358_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6662_ _1863_ _1951_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8401_ _1409_ _3622_ _3354_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ net11 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6898__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5309__I _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6593_ _0844_ _0752_ _1896_ _1898_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8332_ _3552_ _3556_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5544_ _4175_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5570__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7847__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7847__B2 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8263_ as2650.stack\[5\]\[6\] _3241_ _3244_ as2650.stack\[4\]\[6\] _3490_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5475_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7214_ net25 _2475_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8194_ _2781_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7145_ _2414_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _2366_ _2367_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5086__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ as2650.r123\[0\]\[2\] _1373_ _1402_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__A1 _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8575__A2 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7978_ _0403_ _2495_ _3103_ _2480_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _1659_ _1814_ _1811_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8327__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout54 net36 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8878__A3 _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5010__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7838__A1 _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8263__A1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5077__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__I _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6813__A2 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8994__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8566__A2 _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_70 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_81 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_92 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8318__A2 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7609__I _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7829__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4968__I _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5260_ _4069_ _4074_ _4080_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_114_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8884__B _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5191_ _0589_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7057__A2 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8254__A1 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5068__A1 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8950_ _0061_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7901_ _0381_ _3145_ _3146_ _4349_ _2486_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8006__A1 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8881_ _4023_ _4028_ _0555_ _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_13_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7832_ _3014_ _3040_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7763_ _2795_ _3008_ _3012_ _2700_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8124__B _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4975_ _0398_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8309__A2 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__A1 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6714_ _2023_ _2030_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7694_ _2551_ _2362_ _2864_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6645_ _1941_ _1958_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8190__B1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ _1878_ _1885_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6740__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8315_ _3538_ _3520_ _3539_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ _0850_ _0862_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_106_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7296__A2 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8493__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8246_ _3276_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _0839_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8177_ _1023_ _3292_ _3370_ _3070_ _3405_ _0398_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5389_ _4163_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8245__A1 _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7128_ _2403_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__B _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5059__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8085__I _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _0359_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9121__D _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6559__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6534__S _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7429__I _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6333__I _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8720__A2 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8484__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9022__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7039__A2 _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8787__A2 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5412__I _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6798__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9172__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7211__A2 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5222__A1 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4760_ _4353_ _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4576__A3 as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _4273_ _4284_ _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5525__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6722__B2 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6361_ _1668_ _1697_ _1698_ _1213_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8100_ _3132_ _3330_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5312_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9080_ _0177_ clknet_leaf_23_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6292_ _4049_ _0503_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8031_ _1277_ _1511_ _3262_ _3263_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ as2650.addr_buff\[5\] _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5174_ as2650.holding_reg\[0\] _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5322__I _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6789__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7450__A2 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8933_ _0044_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8864_ as2650.psl\[5\] _4008_ _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7815_ _1409_ _2959_ _3063_ _2993_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7202__A2 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8795_ _4367_ _3948_ _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6153__I _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7746_ _2965_ _2880_ _2995_ _2996_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _0356_ _0362_ _0379_ _0382_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6961__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8789__B _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7677_ _2612_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5992__I _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4889_ _0317_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8702__A2 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6628_ _4118_ _1890_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8301__C _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6559_ _4138_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7269__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8466__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8229_ _3426_ _3425_ _3432_ _3433_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8218__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6492__A3 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__B1 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A1 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__B _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A2 _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8154__B1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__A1 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8209__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5691__A1 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__A3 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5930_ as2650.stack\[3\]\[6\] _1310_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _4391_ _1258_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7069__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7600_ _2853_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4812_ _4405_ _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8580_ _4198_ _0438_ _3726_ _3793_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5792_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _2524_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9068__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4743_ as2650.cycle\[10\] _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7462_ _2711_ _2587_ _2714_ _2718_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7499__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8696__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4674_ as2650.ins_reg\[2\] _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8121__C _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6413_ _4364_ _1749_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_128_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7393_ _1718_ _0875_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6171__A2 _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9132_ _0229_ clknet_leaf_33_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8448__A1 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _1666_ _1671_ _1682_ _1670_ _0386_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9063_ _0160_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6275_ _0320_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8014_ as2650.stack\[3\]\[0\] _3246_ _1573_ as2650.stack\[2\]\[0\] _3247_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5226_ _0582_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5052__I _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _0560_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8791__C _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7423__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8620__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5088_ as2650.r123\[3\]\[0\] _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8620__B2 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5434__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4891__I _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8916_ _0027_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8847_ _1139_ _3777_ _3695_ _1534_ _1614_ _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8778_ _2297_ _3931_ _3935_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _2978_ _2979_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7707__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8031__C _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8538__I _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7662__A2 _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4476__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7414__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8273__I _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6925__B2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8222__B _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5137__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8928__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _1392_ _1430_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5011_ _0366_ _0430_ _0431_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6962_ _1209_ _2096_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_81_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8701_ as2650.stack\[5\]\[14\] _3872_ _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5913_ as2650.stack\[3\]\[4\] _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7169__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6893_ _1035_ _2041_ _2097_ _2205_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8632_ as2650.stack\[7\]\[3\] _3835_ _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ as2650.cycle\[0\] _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6916__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7964__I0 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8563_ _0791_ _3777_ _3695_ _2144_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5775_ _0913_ _1156_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_72_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8118__B1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ _2555_ _1672_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4726_ _4319_ _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8669__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8494_ _0420_ _2344_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7971__B _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7445_ _1296_ _1709_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ _4250_ _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7892__A2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7376_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4588_ _4171_ _4180_ _4181_ _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9115_ _0212_ clknet_leaf_38_wb_clk_i as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6327_ _4180_ _1651_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9046_ _0001_ clknet_leaf_14_wb_clk_i as2650.cycle\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7644__A2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6258_ _0606_ _0757_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8841__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5655__A1 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5209_ as2650.psl\[3\] _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _1541_ _1535_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5407__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6606__I _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6080__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8026__C _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__A2 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7955__I0 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6341__I _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7332__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7883__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4697__A2 _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8268__I _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7635__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8832__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8832__B2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7399__A1 _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8217__B _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__I _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6610__A3 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7775__C _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7571__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7347__I _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7571__B2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5560_ _0913_ _0940_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_106_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8887__B _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4511_ as2650.r0\[5\] _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5491_ _0897_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7230_ _4051_ _0340_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7874__A2 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7161_ as2650.r123_2\[0\]\[3\] _2405_ _2435_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6112_ _4253_ _4295_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8823__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7092_ _0533_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ as2650.r123_2\[0\]\[4\] _1375_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8051__A2 _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7994_ _3225_ _3226_ _4057_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _1187_ _2230_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _2181_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7937__I0 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7011__B1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8615_ _1690_ _3738_ _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5827_ _0692_ _1222_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6365__A2 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ as2650.holding_reg\[6\] _4397_ _1159_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8546_ _1678_ _3754_ _3755_ _3761_ _0365_ _0791_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__S1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4709_ _4227_ _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7314__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8477_ _1698_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5689_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7428_ _0542_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5176__I0 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7865__A2 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7359_ _1713_ _2614_ _2617_ _4339_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5505__I as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9124__D _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7617__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9029_ _0140_ clknet_leaf_20_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7720__I _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8290__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8037__B _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8578__B1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A2 _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8042__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5396__B _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A3 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8750__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9129__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9034__D _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7608__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5619__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8281__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6292__A1 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8033__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6044__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7792__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _4253_ _0520_ _1816_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6661_ _1955_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8400_ _3268_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5612_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6592_ _1893_ _1908_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8331_ _3195_ _3532_ _3554_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5543_ _4192_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8262_ as2650.stack\[1\]\[6\] _3242_ _3245_ as2650.stack\[0\]\[6\] _0722_ _3489_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5858__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _4354_ _0387_ _0307_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8193_ _1305_ _3272_ _3421_ _3161_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7144_ _1853_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _2358_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7540__I _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1400_ _1391_ _1372_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6156__I _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6586__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7977_ _3203_ _0433_ _3206_ _3210_ _0334_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6928_ _1144_ _1840_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8304__C _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout55 net32 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7535__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6859_ _2154_ _2155_ _2171_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__9119__D _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5010__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8529_ _1691_ _3745_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5235__I _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6510__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8263__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4824__A2 _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_60 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_71 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_82 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4588__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_93 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8723__B1 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8230__B _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__I _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5190_ _4193_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7057__A3 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8254__A2 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7900_ net52 _0321_ _1519_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8006__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8880_ _1464_ _1475_ _4024_ _4027_ _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_110_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7831_ _2795_ _3075_ _3078_ _2700_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7762_ _2698_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4974_ _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6713_ _2026_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7693_ _2931_ _0461_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7517__A1 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6644_ _1909_ _1937_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8190__A1 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5764__B _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6575_ _1888_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8314_ _0390_ _4073_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5526_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8245_ _3235_ _3471_ _3455_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5457_ _4383_ _0852_ _0858_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_59_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4503__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8176_ _0391_ _2776_ _3404_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5388_ _0778_ _0779_ _0781_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7127_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8245__A2 _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7270__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__C _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5059__A2 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7058_ _2341_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6009_ _1369_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7873__C _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8961__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8484__A2 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6495__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8276__I _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8787__A3 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6798__A2 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7995__A1 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7747__A1 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7211__A3 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5222__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4690_ _4282_ _4283_ _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8172__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7355__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6722__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6360_ _0520_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4733__A1 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _0720_ _0712_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6291_ _0736_ _0738_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_142_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8030_ _1509_ _0338_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6486__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5242_ _0537_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8932_ _0043_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8863_ _0387_ _4010_ _4012_ _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7814_ _2886_ _3058_ _3062_ _4406_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8794_ _4423_ _1249_ _1756_ _1258_ _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5213__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7745_ _2673_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4957_ _4354_ _0298_ _0380_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8789__C _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__A1 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ _2361_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4888_ as2650.cycle\[9\] _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8163__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__I _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _1942_ _1914_ _1943_ _1870_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7265__I _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7910__A1 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A1 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ as2650.holding_reg\[3\] _4377_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6489_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8466__A2 _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8228_ _3445_ _3452_ _3454_ _3455_ _2861_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8218__A2 _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8159_ _3378_ _3357_ _3386_ _3257_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__A1 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5452__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7729__A1 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6401__A1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7884__B _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__A2 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4799__I _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7901__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6704__A2 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7901__B2 _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4715__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A2 _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8209__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__I _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9042__D _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__A4 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _4285_ _1249_ _1260_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8393__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7196__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _4295_ _4255_ _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _1192_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7530_ _2784_ _2785_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4742_ _4335_ _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8145__A1 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7461_ _2715_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4673_ _4266_ _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8696__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _0337_ _0348_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4706__A1 _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _0882_ _0874_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6171__A3 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9131_ _0228_ clknet_leaf_30_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6343_ _1675_ _1681_ _0412_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8448__A2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9062_ _0159_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6274_ _1590_ _1209_ _1594_ _1610_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7120__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5225_ _0613_ _0617_ _0623_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_8013_ _2387_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7959__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5087_ net27 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8620__A2 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6631__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8915_ _0026_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8846_ _1732_ _3171_ _3167_ _3770_ _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8384__A1 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7187__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8777_ as2650.stack\[4\]\[6\] _3932_ _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9012__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5989_ _1268_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7728_ net37 _2932_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7659_ _2808_ _2890_ _4410_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6698__A1 _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9162__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6162__A3 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6870__A1 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4881__B1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8072__B1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8375__A1 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6386__B1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6925__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5728__A3 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4936__A1 _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8127__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8678__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6689__A1 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6249__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8850__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ as2650.cycle\[3\] _0296_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6861__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7789__B _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8063__B1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6961_ _1234_ _2040_ _2270_ _1850_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8700_ _1798_ _3874_ _3881_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5912_ _1271_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8366__A1 _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _2098_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8631_ _2287_ _3834_ _3838_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6377__B1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5843_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6916__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7964__I1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4927__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9185__CLK clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8562_ _1697_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4927__B2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5774_ _0694_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7513_ _2740_ _2768_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6129__B1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4725_ _4315_ _4318_ _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8493_ _3169_ _3710_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7444_ as2650.pc\[3\] _0952_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4656_ _4055_ _4249_ _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5352__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7375_ as2650.pc\[2\] net9 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4587_ _4103_ _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9114_ _0211_ clknet_leaf_29_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6326_ _1090_ _1650_ _0793_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9045_ _0013_ clknet_leaf_13_wb_clk_i as2650.cycle\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6257_ _0995_ _1194_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8841__A2 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ as2650.carry _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6188_ _0674_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5998__I _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ _4082_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6080__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8357__A1 as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8829_ _3344_ _3980_ _3957_ _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6368__B1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7955__I1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4918__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5666__C _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8109__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7580__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7332__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7453__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7096__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8832__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6843__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9058__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8596__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8348__A1 _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__A4 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4761__B _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7571__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4510_ _4103_ _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5490_ _0318_ _0529_ _0324_ _0526_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8520__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4987__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_78_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_78_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7160_ _2153_ _2419_ _2420_ _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5885__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1465_ _0472_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7091_ _2379_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8823__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ as2650.pc\[12\] _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_100_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6834__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7312__B _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8194__I _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5611__I _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8587__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7993_ _3223_ _3222_ _4236_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6944_ _1187_ _2230_ _4092_ _2159_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_54_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6875_ _2184_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7937__I1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7011__A1 as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8614_ _3687_ _1209_ _1589_ _3824_ _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5826_ _0781_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7562__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8545_ _1541_ _1697_ _1698_ _1550_ _3760_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5757_ as2650.holding_reg\[6\] _1057_ _1158_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4708_ as2650.alu_op\[0\] _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8476_ _3687_ _3690_ _3692_ _3693_ _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7314__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8511__A1 _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ _2680_ _2682_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5176__I1 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _4054_ _4228_ _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7865__A3 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5876__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7358_ _2614_ _2616_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _1625_ _1647_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_81_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ _1479_ _0358_ _2548_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6825__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5628__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9028_ _0139_ clknet_leaf_20_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8578__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8578__B2 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4851__A3 _4437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8918__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7250__A1 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8053__B _4448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7002__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6352__I as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8750__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5159__A4 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5564__A1 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7856__A3 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6955__C _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6292__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8569__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7241__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ _4442_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6660_ _1863_ _1951_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5611_ _0988_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6591_ _1894_ _1904_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8330_ _2712_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _0918_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8410__C _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7307__B _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ net9 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8261_ as2650.stack\[3\]\[6\] _3302_ _3303_ as2650.stack\[2\]\[6\] _3488_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4510__I _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7212_ _1517_ _2469_ _2470_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__5858__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8192_ _3221_ _3395_ _3420_ _3391_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7143_ _2404_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4530__A2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__I _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6807__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7074_ as2650.addr_buff\[1\] _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ as2650.r123_2\[0\]\[2\] _1375_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6437__I _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__A3 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A1 _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _1240_ _3207_ _3205_ _3209_ _0465_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _1138_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6858_ _2154_ _2155_ _2171_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7535__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8732__B2 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _0609_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6789_ _4134_ _2048_ _2100_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6900__I _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _4368_ _4218_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8459_ _3537_ _3436_ _3670_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8799__A1 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__B1 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6347__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__I _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4824__A3 _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6791__B _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_61 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_72 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_83 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_127_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A2 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_94 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8723__B2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6966__B _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__A1 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7830_ _2808_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7761_ _3009_ _3010_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7088__I _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6712_ _2024_ _2027_ _2028_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7692_ _2940_ _2942_ _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7517__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6643_ _1938_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8190__A2 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6720__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ _0918_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_wb_clk_i clknet_opt_3_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8313_ _2584_ _4073_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5525_ _0838_ _0847_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8244_ _1674_ _3463_ _3468_ _3470_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ _0854_ _0862_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8647__I _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4503__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8175_ _2767_ _2585_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5387_ _0782_ _0783_ _0790_ _0795_ _0664_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _2402_ _1815_ _2403_ _4343_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5059__A3 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7057_ _2342_ _2343_ _2348_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5071__I _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6008_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7205__A1 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7959_ _3195_ _1674_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8331__B _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8181__A2 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5246__I _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7692__A1 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8557__I _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6495__A2 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7444__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__I _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7995__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8506__B _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7410__B _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4526__S _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5758__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8172__A2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5584__C _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5930__A1 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__I _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A2 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ as2650.psu\[2\] _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6290_ _4449_ _1468_ _0481_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_142_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7683__A1 _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4995__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__A2 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _4230_ _0496_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6238__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7986__A2 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8931_ _0042_ clknet_leaf_32_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5997__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8416__B _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__A3 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8862_ _0306_ _4011_ _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7813_ _1408_ _0377_ _3061_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5749__A1 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5749__B2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8793_ _4235_ _1258_ _1478_ _0429_ _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7744_ _2814_ _2982_ _2994_ _2961_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4956_ _0290_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _2907_ _2924_ _2926_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4972__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4887_ _4351_ _0315_ _0316_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8163__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6174__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ _1873_ _1876_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7910__A2 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ as2650.r123\[0\]\[3\] as2650.r123_2\[0\]\[3\] _4088_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5921__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A2 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _4206_ _0595_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6488_ _4413_ _1802_ _0536_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8227_ _4405_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7674__A1 _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6477__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ as2650.holding_reg\[2\] _0840_ _0843_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_117_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8158_ _1474_ _3369_ _3387_ _0435_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6229__A2 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ as2650.stack\[4\]\[8\] _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8089_ _0785_ _4151_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7977__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9091__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A1 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8840__I _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8154__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__I _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__A1 _4433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7362__B1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4715__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8457__A3 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__B2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7968__A2 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6640__A2 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__I _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__A1 _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8393__A2 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ _4370_ _4403_ _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _1189_ _1190_ _1185_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4741_ _4334_ _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7460_ _2703_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4672_ _4265_ as2650.cycle\[7\] _4266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _1748_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4706__A2 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7391_ _2648_ _2610_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9130_ _0227_ clknet_leaf_33_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6342_ _1676_ _1677_ _1678_ _1680_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_116_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7656__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7315__B _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8197__I _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9061_ _0158_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _1596_ _1611_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5614__I _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8012_ _3244_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5224_ _0626_ _0627_ _0607_ _0628_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8605__B1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _4170_ _0562_ _0563_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_97_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__B1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7959__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5086_ _0433_ _0457_ _0470_ _0505_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8146__B _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6631__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8914_ _0025_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7985__B _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8845_ _3987_ _3980_ _3995_ _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8384__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8951__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8776_ _2295_ _3931_ _3934_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5988_ _1350_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7727_ net38 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4939_ _4047_ _4388_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7276__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7658_ _2905_ _2910_ _2678_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7895__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6698__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6609_ _0601_ _1905_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7589_ _1092_ _1085_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_1_0_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5524__I _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6870__A2 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8072__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8072__B2 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6355__I _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7895__B _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6386__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__B2 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__A4 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__I _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6689__A2 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8063__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8063__B2 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8974__CLK clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7810__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _1228_ _2098_ _1834_ _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6891_ _1017_ _2042_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8366__A2 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8480__I _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8630_ as2650.stack\[7\]\[2\] _3835_ _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6377__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5842_ _4238_ _4288_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6377__B2 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8561_ _3770_ _3775_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5773_ _1169_ _1172_ _1175_ _1176_ _0583_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__4927__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5609__I _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8118__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7512_ _0460_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6129__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4724_ _4249_ _4317_ _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8492_ _1493_ _4308_ _1763_ _4392_ _3709_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_72_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7877__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7443_ _0404_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4655_ _4228_ _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7374_ _2630_ _2631_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _4179_ _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9113_ _0210_ clknet_3_6__leaf_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6325_ _1650_ _1653_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5344__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9044_ _0012_ clknet_leaf_21_wb_clk_i as2650.cycle\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6256_ _1160_ _1163_ _1065_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6301__A1 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _0608_ _0612_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6187_ _0778_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5138_ _4449_ _0493_ _0546_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A3 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8357__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8828_ _2473_ _1752_ _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6368__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6368__B2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__A2 _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8759_ _1238_ _3906_ _3922_ _3923_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8109__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A2 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7868__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5254__I _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8293__A1 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7096__A2 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8045__A1 _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8514__B _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7859__A1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8520__A2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6531__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _4060_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8284__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _2377_ _2378_ _2359_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9002__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8475__I _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _1370_ _1414_ _1415_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5893__I0 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ _3222_ _3223_ _3224_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9152__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6943_ _2252_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5270__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _2185_ _2160_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8613_ _3734_ _1234_ _3823_ _3687_ _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5825_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5339__I _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8544_ _0815_ _3350_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5756_ as2650.holding_reg\[6\] _1158_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ _4294_ _4300_ _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8475_ _2943_ _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7554__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5687_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7426_ _2680_ _2682_ _2614_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4638_ _4072_ _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6522__A1 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7357_ _2569_ _2615_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4569_ _4160_ _4077_ _4161_ _4070_ _4162_ _4067_ _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5074__I _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6308_ _1628_ _1631_ _1637_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7288_ _4442_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9027_ _0138_ clknet_leaf_73_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _1577_ _1404_ _1582_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4836__A1 _4424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8578__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A4 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8334__B _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8750__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8502__A2 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6513__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9025__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8266__B2 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9175__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8228__C _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8569__A2 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7241__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5610_ _0780_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6590_ _0876_ _1906_ _1901_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5541_ _0944_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ _2497_ _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5307__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ _4207_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7211_ _2473_ _4353_ _0291_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8191_ _3410_ _3419_ _2731_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5858__A3 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8257__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7142_ _2403_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4530__A3 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6807__A2 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7073_ _1713_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5622__I _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8138__C _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _1399_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__C _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A2 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ _0300_ _2498_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _1831_ _2222_ _2237_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5794__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _2168_ _2170_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_74_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5069__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8732__A2 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5808_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6743__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _4214_ _1814_ _2101_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8527_ _1677_ _1695_ _3742_ _3743_ _3310_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5739_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__B _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__I _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8496__A1 _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8458_ _3672_ _3676_ _3232_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7409_ _2551_ _2639_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5849__A3 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8389_ _3367_ _3610_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__A4 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8799__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__A1 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4809__B2 _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__A3 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6363__I _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_62 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_73 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_84 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6982__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4588__A3 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_95 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8184__B1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8723__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6734__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__A2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8487__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8239__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__A2 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7214__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8411__A1 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7760_ net38 net37 _2932_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _4295_ _4261_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5776__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _4117_ _1861_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7691_ _2574_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _1941_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5528__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8421__C _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5617__I _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8312_ _3512_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8478__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8243_ _3027_ _3469_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5455_ _0854_ _0862_ _0621_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__A1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8174_ _2596_ _3394_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5700__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ _0791_ _0794_ _0783_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7053__B _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7125_ _1131_ _1828_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7056_ _4323_ _0516_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5464__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ as2650.r123\[0\]\[0\] _1373_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7756__A3 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7958_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6909_ _1078_ _2059_ _2219_ _2220_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7889_ _3108_ _3131_ _3134_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8331__C _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6192__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8985__D _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7742__I _4440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5262__I _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7444__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8641__A1 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__I _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5758__A2 _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6955__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7917__I _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6707__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7380__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5930__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _4193_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7683__A2 _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8880__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _4389_ _4299_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7435__A2 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8483__I _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8930_ _0041_ clknet_leaf_36_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5997__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7199__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8861_ _0931_ _0996_ _1008_ _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7099__I _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4516__I _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7812_ _2553_ _3052_ _3060_ _2989_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8792_ _3943_ _3944_ _3945_ _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _2965_ _2959_ _2992_ _2993_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4955_ _4445_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__I _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7674_ _2759_ _2925_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4886_ _4337_ _0296_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7048__B _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6625_ _4117_ _1874_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7371__A1 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6174__A2 _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5347__I _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7910__A3 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _4117_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5921__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5507_ _0856_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7123__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6487_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _3260_ _3425_ _3453_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _0845_ _0587_ _4395_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8871__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8157_ _2472_ _3372_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5369_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5082__I _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _2391_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8088_ _1716_ _4135_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7039_ _0443_ _4275_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A2 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__A1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6165__A2 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7362__B2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7472__I _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8862__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8614__A1 _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6928__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__B2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ _4332_ _4333_ _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4671_ _4264_ _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5167__I _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ _1689_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9109__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7390_ _0786_ _0802_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5903__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4706__A3 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6341_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9060_ _0157_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6272_ _0608_ _0758_ _0854_ _1600_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5667__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8011_ _3243_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6864__B1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ _0629_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8605__A1 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5154_ _4297_ _0473_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8427__B _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4890__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6726__I _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5085_ _0500_ _0504_ _4363_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8913_ _0024_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8369__B1 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A2 _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6919__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8844_ _1630_ _3991_ _3994_ _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7592__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A2 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5987_ _1331_ _1360_ _1365_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8775_ as2650.stack\[4\]\[5\] _3932_ _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6461__I _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7726_ _2566_ _2974_ _2976_ _2744_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4938_ _4341_ _4304_ _4380_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7344__A1 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7657_ _2562_ _2908_ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6608_ _0777_ _1906_ _1922_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7895__A2 _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7588_ _1093_ _1085_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6539_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7292__I _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8844__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5658__A1 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8209_ _0533_ _2334_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9189_ _0286_ clknet_leaf_43_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6572__S _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7895__C _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6386__A2 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6371__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7335__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5715__I as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8063__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6074__A1 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7810__A2 _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8761__I _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _1303_ _1273_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6890_ _0880_ _2045_ _2099_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_46_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8366__A3 _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5841_ _0720_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6377__A2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _1162_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8560_ _3771_ _3773_ _3774_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__A3 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7511_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4723_ _4268_ _4316_ _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8491_ _4299_ _4315_ _4385_ _0572_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6129__A2 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7442_ _2678_ _2695_ _2697_ _2698_ _4410_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7877__A2 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4654_ _4232_ _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9081__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7373_ net30 _2540_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4585_ _4173_ _4175_ _4177_ _4178_ _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_116_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9112_ _0209_ clknet_leaf_27_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _1654_ _4370_ _1655_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8826__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9043_ _0011_ clknet_leaf_15_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _1009_ _1078_ _1177_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_143_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6301__A2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _0615_ _4251_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6186_ _1530_ _1537_ _1539_ _1508_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ _0518_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_85_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5068_ _4398_ _0478_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__B1 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8827_ _3979_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__A2 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__I _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8758_ _3892_ _2276_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _0386_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8689_ _1781_ _3873_ _3875_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8817__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6828__B1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7750__I _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6056__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5803__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8348__A3 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A1 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7925__I _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__B1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7859__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A1 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5445__I _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6531__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8808__A1 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8284__A2 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ as2650.stack\[1\]\[11\] _1397_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5893__I1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7991_ _1217_ _4188_ _4220_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_81_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _2229_ _2231_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5270__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_16_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7547__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ _2128_ _2158_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8612_ _3765_ _1228_ _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ _0672_ _0959_ _1224_ _1032_ _1226_ _0871_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_5755_ _4181_ _4396_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8543_ _3756_ _3757_ _1700_ _3758_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4781__A1 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _4296_ _4298_ _4299_ _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5686_ net1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8474_ _3691_ _0638_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7425_ _2641_ _2642_ _2681_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4637_ _4226_ _4230_ _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6522__A2 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7356_ _1712_ _0806_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4568_ as2650.r123\[1\]\[0\] as2650.r123\[0\]\[0\] as2650.r123_2\[1\]\[0\] as2650.r123_2\[0\]\[0\]
+ as2650.ins_reg\[0\] _4062_ _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _0490_ _1641_ _1642_ _0302_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_7287_ _2538_ _2539_ _2543_ _2546_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _4059_ _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9026_ _0137_ clknet_leaf_74_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6238_ as2650.stack\[3\]\[10\] _1580_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__A2 _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _0385_ _4420_ _1521_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_44_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6038__A1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7786__A1 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8988__D _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7745__I _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6761__A2 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7710__A1 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7710__B2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5721__B1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7480__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6277__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4827__A2 _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__A1 as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8525__B _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6201__A1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5540_ _0945_ _0648_ _0946_ _0649_ _4134_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_121_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ _0667_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5175__I _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7210_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8190_ _3378_ _3395_ _3415_ _3257_ _3418_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7141_ _2418_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8257__A2 _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _2329_ _2360_ _2364_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6023_ as2650.pc\[10\] _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7768__A1 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _1655_ _1722_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6925_ as2650.r123_2\[2\]\[5\] _2112_ _2236_ _2142_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _2122_ _2136_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout47 net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5794__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ _1187_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8987__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7940__A1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _2046_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8526_ _1534_ _1697_ _1698_ _0950_ _1639_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5738_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8496__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8457_ _0656_ _3463_ _3162_ _3675_ _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5669_ _0995_ _0999_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7408_ _2335_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8388_ _2374_ _2553_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7339_ _1499_ _2597_ _1288_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__I _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6259__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8329__C _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8799__A3 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__A2 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9009_ _0120_ clknet_leaf_78_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A2 _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_63 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_74 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_85 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_96 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8184__B2 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8080__B _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7931__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8487__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__A1 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9142__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8239__A2 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7998__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _4443_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _4127_ _1857_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4984__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7690_ _2607_ _2941_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8175__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _1946_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7922__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7318__C _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ as2650.r123\[0\]\[2\] as2650.r123_2\[0\]\[2\] _4108_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8311_ _3533_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5523_ _0620_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8478__A2 _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8242_ _3464_ _3467_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5454_ _0765_ _0860_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_117_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5161__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6729__I _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8173_ _2864_ _3400_ _3401_ _2354_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5385_ _0428_ _0493_ _0547_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_82_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7124_ _0573_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7055_ _2344_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6006_ _1374_ _1377_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5464__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_86_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6413__A1 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7957_ _2407_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6908_ _1086_ _1826_ _2059_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7888_ _0385_ _3132_ _2486_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _0940_ _2096_ _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7295__I _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5519__A3 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__I _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7913__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4727__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8509_ _3726_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7244__B _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5543__I _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7898__C _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6374__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5207__A2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6404__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6307__C _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6955__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A1 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7904__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6707__A2 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5718__I _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A1 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7933__I _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6891__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5170_ _0567_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8860_ _3802_ _4009_ _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8396__A1 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7199__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7811_ _3049_ _4431_ _2721_ _3059_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8791_ _0449_ _1471_ _0428_ _0677_ _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4957__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7742_ _4440_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4954_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9188__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7673_ _2584_ _1227_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8699__A2 _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _0313_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4532__I _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _1939_ _1892_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7048__C _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6555_ _1871_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ _0567_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7123__A2 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6486_ _0524_ _4374_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8225_ _2407_ _3435_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5437_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8871__A2 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8608__C1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8156_ _0831_ _3383_ _3384_ _3385_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8674__I _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8087_ _2664_ _3317_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5299_ _0707_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8623__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8607__C _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7038_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8387__A1 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8989_ _0100_ clknet_leaf_9_wb_clk_i as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8139__A1 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__A2 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7114__A2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8862__A2 _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__I _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8075__B1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8614__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__B1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6928__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7050__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4939__A1 _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8252__C _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4670_ _4263_ _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5364__A1 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _0953_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8302__A1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7105__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6271_ _1590_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8853__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5222_ _4390_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8010_ _0699_ _0701_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6864__B2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _4282_ _0492_ _0542_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8605__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5911__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _4236_ _4257_ _4446_ _0503_ _4312_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8912_ _0023_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8369__A1 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8369__B2 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8843_ _3772_ _0479_ _3992_ _3993_ _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6919__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5786__C _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8774_ _2291_ _3931_ _3933_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ as2650.stack\[1\]\[7\] _1361_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8162__C _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6395__A3 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7725_ _2971_ _2975_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ _0298_ _0358_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _2903_ _2564_ _2612_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4868_ _4428_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7344__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8541__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _0601_ _1923_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5355__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7587_ _2840_ _1153_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _4079_ _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6538_ _1729_ _1829_ _1854_ _0322_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6469_ _1789_ _1786_ _1791_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8208_ _0737_ _0376_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5658__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9188_ _0285_ clknet_leaf_44_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8618__B _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7522__B _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8139_ _2710_ _3356_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6607__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7804__B1 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8780__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8532__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8800__C _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5346__B2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__A1 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6827__I _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8366__A4 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ _1182_ _0983_ _1239_ _1242_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _0770_ _1165_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5178__I _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ as2650.pc\[4\] _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _4052_ _4157_ _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8490_ _2993_ _1839_ _1691_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8523__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7441_ _2620_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4653_ _4242_ _4246_ _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7877__A3 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__B _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ net31 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ _4129_ _4132_ _4136_ _4141_ _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_128_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9111_ _0208_ clknet_leaf_27_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ _0476_ _1659_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9042_ _0010_ clknet_leaf_40_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6254_ _0638_ _0940_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ net42 _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5641__I _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _4438_ _0447_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7262__A1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _4384_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7996__C _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__B1 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8826_ _1689_ _3978_ _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8757_ as2650.r123\[2\]\[7\] _3912_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5969_ _1353_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4918__A4 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7708_ _1381_ _2534_ _2958_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8688_ as2650.stack\[5\]\[8\] _3874_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8514__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5328__A1 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7639_ _2550_ _2384_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4720__I _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8278__B1 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8817__A2 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6828__A1 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__B2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7252__B _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7253__A1 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4606__A3 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7005__A1 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8753__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A3 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8505__A1 _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8530__C _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7859__A3 _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4542__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7492__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8772__I _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7990_ _1275_ _0429_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _2227_ _2228_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__A3 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6872_ _2128_ _2158_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6225__C _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8611_ _3731_ _3821_ _3822_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5823_ _4081_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8542_ _2005_ _0572_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5754_ _4103_ _0541_ _1157_ _4378_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_56_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4705_ _4233_ _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4781__A2 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8473_ _3686_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5685_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8012__I _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7424_ _1717_ _0893_ _0895_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4636_ _4229_ _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7355_ _0542_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5730__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _4062_ _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _1473_ _1644_ _1515_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7286_ _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4498_ _4091_ _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7483__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6467__I _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9025_ _0136_ clknet_leaf_71_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6286__A2 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _1577_ _1396_ _1581_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5494__B1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6168_ _4416_ _0315_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ as2650.cycle\[5\] as2650.cycle\[4\] _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6099_ as2650.r123_2\[3\]\[6\] _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8735__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5549__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8809_ _0733_ _0973_ _3962_ _3195_ _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8350__C _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5546__I _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6277__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7226__A1 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6029__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__B1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__B _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9071__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7529__A2 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _0688_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7140_ as2650.r123_2\[0\]\[0\] _2405_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6268__A2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ _2362_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5191__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6022_ _1370_ _1396_ _1398_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7217__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8435__C _4424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7973_ _2510_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6924_ _2223_ _2225_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _2124_ _2135_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6786_ _0882_ _2049_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5400__B1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7940__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8525_ _3737_ _3741_ _1701_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5737_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8456_ as2650.pc\[14\] _3674_ _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5668_ _0986_ _0991_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7407_ _2664_ _0305_ _2533_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4619_ _4156_ _4166_ _4195_ _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8387_ _1408_ _3608_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5599_ _0615_ _0496_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7338_ _2596_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6197__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7456__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6259__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7269_ _1252_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8799__A4 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9008_ _0119_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9094__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A1 _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8345__C _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_75 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_86 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8931__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8184__A2 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7931__A2 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5942__A1 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7695__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7705__B _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_1_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7998__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4681__A1 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4970_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8271__B _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8175__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _1947_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_75_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7922__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4736__A2 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _1880_ _1886_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5186__I as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8310_ _4425_ _3473_ _3534_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5522_ _0925_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7686__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8241_ _3464_ _3467_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _0750_ _0756_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8172_ _1672_ _2335_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5161__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5384_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7123_ _1800_ _2393_ _2401_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _0404_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _1381_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4672__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8954__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6413__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_71_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_71_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7956_ _3193_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6907_ _2097_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7887_ _1258_ _0430_ _0679_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _0948_ _2040_ _2151_ _2057_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7509__C _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7913__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _1968_ _1860_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8508_ _1628_ _3711_ _3716_ _3725_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_109_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8439_ _3650_ _3651_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7244__C _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8075__C _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8157__A2 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A2 _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7668__A1 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5734__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8617__B1 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8977__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[33] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7810_ _2550_ _3044_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8790_ _2471_ _0388_ _2336_ _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _2886_ _2986_ _2991_ _4406_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4957__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4953_ _4420_ _0366_ _0374_ _0377_ _4257_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7672_ _0390_ _1227_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6159__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4884_ _4332_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6623_ _1878_ _1885_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ as2650.r123\[0\]\[1\] as2650.r123_2\[0\]\[1\] _4088_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7659__A1 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5505_ as2650.r123\[0\]\[3\] _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6485_ _0337_ _4245_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8320__A2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8224_ _3281_ _3425_ _3451_ _2548_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _4139_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4568__S1 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8155_ as2650.stack\[1\]\[3\] _2456_ _3254_ as2650.stack\[0\]\[3\] _0825_ _3385_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8608__B1 _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5367_ _0752_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8608__C2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8084__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8086_ _2582_ _1275_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5298_ as2650.psu\[1\] _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7831__A1 _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7037_ _0562_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A1 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6398__B2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9132__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8988_ _0099_ clknet_leaf_9_wb_clk_i as2650.alu_op\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7939_ _1545_ _1499_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7898__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7255__B _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8847__B1 _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5125__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6322__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6625__A2 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__I as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__B2 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7050__A2 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4939__A2 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4633__I _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7889__A1 _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6936__I0 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7105__A3 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6270_ _1607_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6313__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _4303_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6864__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7813__A1 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4808__I _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4627__A1 _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9155__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8911_ _0022_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8842_ _1212_ _2472_ _1626_ _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8773_ as2650.stack\[4\]\[4\] _3932_ _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5985_ _1325_ _1360_ _1364_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4543__I _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ _2972_ _2920_ _2921_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4936_ _4400_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ _0391_ _1228_ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4867_ _4365_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6606_ _1898_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7586_ _1140_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4798_ _4303_ _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_119_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6537_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5374__I _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ as2650.stack\[6\]\[9\] _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8207_ _2586_ _2819_ _3434_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ as2650.stack\[3\]\[9\] _0714_ _0704_ as2650.stack\[1\]\[9\] _0828_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9187_ _0284_ clknet_leaf_67_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ _1210_ _1524_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4866__A1 _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8057__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8138_ _2864_ _3366_ _3367_ _2354_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7804__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6607__A2 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7804__B2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8069_ _4362_ _3275_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__A1 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8353__C _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__I _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6791__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5284__I _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8296__A1 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__A2 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9178__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8048__A1 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8599__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4628__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4609__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8544__B _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _0625_ _1173_ _1163_ _1005_ _0914_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_72_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _4252_ _4239_ _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7440_ net55 _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _4245_ _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6511__C _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7371_ _2581_ _2627_ _2628_ _2629_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _4147_ _4153_ _4176_ _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_122_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9110_ _0207_ clknet_leaf_24_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6322_ _1660_ _1658_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__B _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9041_ _0009_ clknet_leaf_13_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6253_ _0775_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4848__A1 _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _4389_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6184_ _1529_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _0368_ _0302_ _0519_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _4387_ _4248_ _0473_ _4382_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_84_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8173__C _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__A1 _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8211__B2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8825_ _1349_ _3975_ _3977_ _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8756_ _1179_ _3906_ _3921_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4919_ as2650.cycle\[7\] _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7707_ _2728_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5899_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8687_ _3872_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7638_ _2720_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5328__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6525__A1 _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7569_ _2722_ _2811_ _2823_ _0440_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8278__A1 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9239_ net48 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7252__C _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8825__I0 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7253__A2 _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7759__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7005__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__I _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6764__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4911__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A3 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7492__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A3 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7244__A2 _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5255__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6573__I _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _2232_ _2233_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _2182_ _2183_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5189__I _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ _4179_ _4103_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8610_ _1319_ _3750_ _0351_ _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6755__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ _4100_ _0541_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8541_ _1350_ _3698_ _0573_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5917__I _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4821__I _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _4297_ _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6507__A1 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8472_ _3688_ _0660_ _3689_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5684_ _4104_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7423_ _1710_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _4227_ _4228_ _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7180__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _1713_ _2561_ _2609_ _2611_ _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4566_ _4159_ _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4977__B _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5730__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _1643_ _0731_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7285_ _2471_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4497_ _4090_ _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9024_ _0135_ clknet_leaf_5_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6236_ as2650.stack\[3\]\[9\] _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7483__A2 _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6167_ _1518_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7235__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5118_ _4347_ _4333_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_111_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _1455_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8735__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8808_ _3959_ _3960_ _3961_ _0733_ _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7528__B _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8739_ _0696_ _3906_ _3910_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6432__B _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8499__A1 _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7171__A1 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5562__I _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6277__A3 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8671__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7226__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__B2 _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6434__B1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6985__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__C _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8113__I _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4920__B1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9091__D _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5472__I _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7070_ _2358_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8662__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5476__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ as2650.stack\[1\]\[9\] _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7870__C1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8414__A1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7217__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4816__I _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6976__A1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7972_ _3111_ _3205_ net4 _2510_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6923_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8717__A2 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _2157_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5805_ _0914_ _1185_ _1198_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6785_ _1817_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5400__B2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5736_ net2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8524_ _1922_ _0503_ _3740_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7153__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5667_ _0855_ _1066_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8455_ _3441_ _3673_ _1756_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7862__I _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8350__B1 _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7406_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4618_ _4207_ _4211_ _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8386_ _2999_ _3563_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ _0616_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5703__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7337_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4549_ _4137_ _4142_ _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5382__I _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7268_ _4401_ _2478_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7456__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6219_ net21 _1559_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7811__B _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9007_ _0118_ clknet_leaf_78_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7199_ _2459_ _1414_ _2465_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8405__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A2 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A1 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5050__C _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_65 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7392__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__I _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5942__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7695__A2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7705__C _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8892__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8644__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8108__I _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6186__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7383__A1 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5467__I _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__A3 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _1881_ _1883_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4736__A3 _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _0770_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7135__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8240_ _3465_ _3448_ _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _0606_ _0619_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8883__A1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5697__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8171_ _1022_ _4120_ _3399_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5383_ _4419_ _0447_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7122_ as2650.stack\[4\]\[14\] _2391_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5449__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7053_ _0329_ _2345_ _0323_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _0555_ _1267_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4672__A2 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8018__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7955_ _1503_ _1056_ _3186_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5621__A1 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6906_ _2212_ _2098_ _2217_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7886_ _0360_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8020__C1 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _0962_ _2041_ _1834_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7374__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4727__A3 _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6768_ _2080_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7806__B _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8507_ _1642_ _3717_ _3721_ _3724_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7126__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5719_ _1122_ _0818_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6699_ _2014_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_109_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8438_ _3653_ _3655_ _3656_ _3657_ _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8874__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9061__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8369_ _4425_ _3588_ _3590_ _3591_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__I _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8356__C _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A2 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4456__I _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7601__A2 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5287__I _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7668__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5143__A3 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8880__A4 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8617__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8617__B2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8547__B _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7451__B _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__S _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8093__A2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__I _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5851__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 io_in[34] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7677__I _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7740_ _2965_ _0377_ _2990_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4952_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4957__A3 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7671_ _2361_ _2922_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4883_ as2650.cycle\[1\] _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7356__A1 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6159__A2 _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6622_ _1878_ _1885_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _4105_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5504_ _0836_ _0578_ _0911_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4590__A1 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__C _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7659__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6484_ _1800_ _1787_ _1801_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8856__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8223_ _2723_ _3449_ _3450_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5435_ _4137_ _4142_ _0599_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8608__A1 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _0762_ _0769_ _0774_ _0750_ _0583_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_8154_ as2650.stack\[3\]\[3\] _3302_ _1574_ as2650.stack\[2\]\[3\] _3384_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8608__B2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7105_ _1243_ _2389_ _1782_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8085_ _2731_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8084__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7036_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7831__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7595__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8987_ _0098_ clknet_leaf_1_wb_clk_i as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _3179_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7869_ _2507_ _3100_ _3115_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7898__A2 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__C _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8847__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8847__B2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6322__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8075__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6086__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4914__I _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7050__A3 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7165__C _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4572__A1 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8838__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8944__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6313__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5220_ _0370_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5151_ _4356_ _4344_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8066__A2 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7813__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5082_ _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4627__A2 _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8910_ _0021_ clknet_leaf_76_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7026__B1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8841_ _3169_ _3952_ _0574_ _1636_ _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8772_ _3924_ _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ as2650.stack\[1\]\[6\] _1361_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7723_ _2971_ _2973_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7329__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7654_ _2834_ _2833_ _2835_ _2906_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _4429_ _4444_ _0297_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6605_ _1896_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7585_ _2760_ _2837_ _2838_ _2693_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4797_ _4390_ _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8829__A1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6536_ _0740_ _1812_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7501__A1 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6467_ _1784_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8206_ _1314_ _4415_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5418_ _0709_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9186_ _0283_ clknet_leaf_44_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6398_ _1731_ _1734_ _1735_ _1690_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4866__A2 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8057__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8137_ _1680_ _2863_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5349_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7804__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8068_ _3175_ _3290_ _0414_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _2301_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7017__B1 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7568__A1 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6154__C _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8967__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7740__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8296__A2 _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8809__C _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8048__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__I as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6059__A1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__B _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4644__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8116__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4720_ _4313_ _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _4243_ _4244_ _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7731__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5475__I _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7370_ _1507_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _4163_ _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ as2650.psl\[6\] _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6298__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9040_ _0008_ clknet_3_2__leaf_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6252_ _0839_ _0865_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_143_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _0608_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_115_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6183_ _0698_ _1533_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5134_ _0317_ _0528_ _0538_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _0475_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4554__I _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8824_ _3426_ _3976_ _3957_ _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8211__A2 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8755_ _3900_ _2261_ _3909_ as2650.r123\[2\]\[6\] _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5967_ _1346_ _1347_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7970__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7706_ _2948_ _2957_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4918_ _0309_ _4282_ as2650.cycle\[12\] _4270_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_40_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8686_ _3872_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5898_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7637_ net54 _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7722__A1 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4849_ _4441_ _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7568_ _2809_ _2601_ _2723_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8278__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ _1820_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7499_ _0953_ _0961_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6289__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9238_ net48 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4729__I _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9169_ _0266_ clknet_leaf_4_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8825__I1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7253__A3 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8450__A2 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9179__D _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8738__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6764__A2 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4775__A1 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5295__I _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9145__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8269__A2 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5255__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6870_ _4076_ _1864_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ _0671_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8540_ as2650.overflow _3701_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5752_ _1151_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ _4053_ _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8471_ _2762_ _0651_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7704__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4518__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7422_ _0944_ _0947_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4634_ as2650.alu_op\[2\] _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7180__A2 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__B _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ _2345_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4565_ as2650.r0\[0\] _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6304_ _1265_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7284_ _4441_ _0397_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4496_ _4089_ _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9023_ _0134_ clknet_leaf_74_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6235_ _1575_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8680__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4541__I1 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _1513_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5117_ _4045_ _4261_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6097_ as2650.r123_2\[3\]\[5\] _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _4259_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9018__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__A1 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8807_ _0877_ _3959_ _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6746__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6999_ _2299_ _2292_ _2300_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4757__A1 _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8738_ _3900_ _2036_ _3909_ as2650.r123\[2\]\[0\] _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8499__A2 _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8669_ _2285_ _3859_ _3862_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5706__B1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A1 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__I _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__I _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5485__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8375__B _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7226__A3 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6434__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__B2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8187__A1 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4920__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8111__A1 _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8662__A2 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _1368_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7901__C _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7870__B1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__C2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7217__A3 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7971_ _3203_ _0394_ _3204_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6922_ _2232_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8178__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ _2164_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _0930_ _1204_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6784_ _1821_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8523_ _0702_ _3738_ _0574_ _3739_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5735_ _0672_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8454_ _3671_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5666_ _0626_ _1069_ _1070_ _0632_ _0582_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8350__A1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8350__B2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ as2650.pc\[2\] _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4617_ _4192_ _4209_ _4210_ _4196_ _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8385_ _2713_ _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5597_ _0995_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7336_ _4324_ _4313_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4548_ _4141_ _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8102__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8653__A2 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7267_ _1277_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4479_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _4064_ _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9006_ _0117_ clknet_leaf_78_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ _1319_ _1555_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7198_ as2650.stack\[2\]\[11\] _2462_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6494__I _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ as2650.psu\[5\] _1491_ _1498_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6416__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A2 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_as2650_88 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7916__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A4 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4742__I _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7392__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8892__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A1 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8644__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__A3 _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7907__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__I _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8580__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7922__A4 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4736__A4 _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _0853_ _0926_ _4383_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7135__A2 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__I _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _0586_ _0592_ _0593_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6894__A1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5697__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8170_ _3398_ _3365_ _3361_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5382_ _4144_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7121_ _1798_ _2393_ _2400_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5449__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7052_ _4265_ _4337_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8399__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7071__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7954_ _3192_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6905_ _1087_ _2044_ _1835_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7885_ _0432_ _2487_ _3127_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_35_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8020__B1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6836_ _2043_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5385__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ as2650.r0\[4\] _1857_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _2344_ _3723_ _1528_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5718_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8323__A1 _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6698_ _4150_ _1973_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7126__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8323__B2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6489__I _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8437_ _2374_ _2378_ _3590_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5649_ as2650.r123\[0\]\[5\] _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_80_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8368_ _2371_ _3589_ _2354_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ _2527_ _2530_ _2578_ _0458_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8299_ _3512_ _3502_ _3519_ _3238_ _3524_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_49_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5860__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8372__C _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6173__B _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9187__D _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8314__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7117__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8865__A2 _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8617__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4647__I _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5851__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput7 io_in[5] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4957__A4 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7670_ _2920_ _2921_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ _0308_ _0312_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7356__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6621_ _1888_ _1891_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_75_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6552_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5503_ _0579_ _0901_ _0910_ _0577_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6483_ as2650.stack\[6\]\[14\] _1785_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8856__A2 _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8222_ _1095_ _2552_ _3234_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6867__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5434_ as2650.holding_reg\[2\] _0840_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8153_ as2650.stack\[7\]\[3\] _2389_ _3380_ as2650.stack\[4\]\[3\] _3382_ _3383_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5365_ _0770_ _0758_ _0773_ _0636_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5941__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8084_ _1288_ _3272_ _3315_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5296_ as2650.psu\[0\] _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7035_ _1708_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A2 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7044__A1 _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8986_ _0097_ clknet_leaf_3_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8192__C _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8792__A1 _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7937_ _3178_ as2650.holding_reg\[1\] _3166_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7868_ _3101_ _3114_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8544__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _2127_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7799_ _2566_ _3046_ _3047_ _2744_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8847__A2 _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6307__B1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7108__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6012__I as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5530__A1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__I as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8783__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5597__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__I as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7889__A3 _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__A2 _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8838__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8558__B _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__B _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _0517_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5081_ _4297_ _4094_ _0473_ _4382_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_99_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7026__A1 as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7026__B2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8840_ _3990_ _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5037__B1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8774__A1 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8771_ _3924_ _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9051__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _1317_ _1360_ _1363_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7722_ _2907_ _2924_ _2926_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_75_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4934_ _4280_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_19_wb_clk_i clknet_opt_2_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7329__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8526__B2 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7653_ _2898_ _1138_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4865_ as2650.cycle\[12\] _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5936__I _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8312__I _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6604_ _1918_ _1919_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _1673_ _2760_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4796_ _4389_ _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8829__A2 _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _1395_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7501__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8205_ _3257_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5512__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ as2650.stack\[5\]\[9\] _0824_ _0726_ as2650.stack\[4\]\[9\] _0825_ _0826_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_9185_ _0282_ clknet_3_7__leaf_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6397_ _1692_ _1476_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8136_ _3363_ _3365_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5348_ _0750_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8067_ _3278_ _3280_ _3275_ _3282_ _3298_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5279_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _2153_ _2302_ _2315_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7568__A2 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5579__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8969_ _0080_ clknet_leaf_15_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6240__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7547__B _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7740__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8378__B _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6551__I0 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7008__A1 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7301__I _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8756__A1 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__C _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8841__B _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8508__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8911__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4650_ net5 _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7731__A2 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 io_in[8] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5742__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _4174_ _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6320_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6251_ _0615_ _4392_ _4450_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_131_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4848__A3 _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ _1534_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7247__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5133_ _4338_ _0542_ _0530_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7920__B _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7798__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _0479_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8307__I _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__I _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8823_ _1499_ _1677_ _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8754_ _3919_ _3920_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _1349_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7970__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7705_ _2931_ _0393_ _2714_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4917_ _0335_ _0344_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8685_ _3871_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5981__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ as2650.pc\[3\] _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_90_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4570__I _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7636_ net35 net34 _2810_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4848_ _4296_ _4278_ _4240_ _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7567_ _2821_ _1502_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4779_ _4372_ _4086_ _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6518_ _1805_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7498_ _2736_ _0961_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9237_ net47 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7486__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6497__I _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6289__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ as2650.stack\[0\]\[11\] _1774_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9168_ _0265_ clknet_leaf_78_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9097__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8435__B1 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8119_ _3345_ _3346_ _3348_ _3349_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9099_ _0196_ clknet_leaf_82_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7253__A4 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__I _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8934__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__B1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A2 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__I as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7992__S _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__A2 _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7477__A1 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7740__B _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4655__I _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5820_ _4181_ _1079_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _0643_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4295_ _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8470_ _2566_ _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5682_ _4106_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7704__A2 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6507__A3 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8901__A1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7421_ _0324_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4518__A2 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _4054_ _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7352_ _2560_ _2610_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _4052_ _4054_ as2650.alu_op\[2\] _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_116_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7468__A1 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _0369_ _0363_ _0364_ _0372_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7283_ _2541_ _2542_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4495_ as2650.r123\[0\]\[6\] as2650.r123_2\[0\]\[6\] _4088_ _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9022_ _0133_ clknet_leaf_5_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6110__I _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6234_ _1577_ _1386_ _1579_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6691__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6165_ _4433_ _4344_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8465__C _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5116_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _1454_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7640__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6443__A2 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4565__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8957__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5047_ _0436_ _0464_ _0465_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_34_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_84_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8806_ _1350_ _1574_ _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6998_ as2650.stack\[5\]\[7\] _2293_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4757__A2 _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8737_ _3908_ _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5949_ _1300_ _1334_ _1339_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8668_ as2650.stack\[6\]\[1\] _3860_ _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8499__A3 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7619_ _1322_ _2533_ _0320_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8599_ _3765_ _1154_ _3691_ _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5345__B _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__I _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__A1 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7560__B _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__B _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6434__A2 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5642__B1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__I0 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__A2 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9112__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4920__A2 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__B2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__C _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A1 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7622__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7970_ _0472_ _1694_ _1495_ _1654_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6921_ _2161_ _2163_ _2188_ _2189_ _2180_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _2127_ _2133_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6189__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _0628_ _1195_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4739__A2 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _1806_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8522_ as2650.psl\[1\] _3698_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5734_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7689__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8453_ _1429_ _3473_ _3671_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5665_ _1062_ _1064_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7404_ _1694_ _2660_ _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8350__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _4157_ _4158_ _4165_ _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8384_ _1408_ _2538_ _3605_ _4049_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6361__A1 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ _0849_ _0937_ _0926_ _0922_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6361__B2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7335_ _2546_ _2591_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _4139_ _4077_ _4140_ _4067_ _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_116_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8102__A2 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7266_ _2525_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4478_ _4071_ _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9005_ _0116_ clknet_leaf_79_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7861__A1 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ _1090_ _1556_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7197_ _2459_ _1404_ _2464_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _1499_ _1502_ _1492_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_85_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7613__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6416__A2 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ as2650.stack\[0\]\[4\] _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_56 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_57_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7916__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__I _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4902__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7852__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4933__I _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8565__C1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5918__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8580__A2 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8140__I _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5450_ _0632_ _0853_ _0854_ _0628_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9008__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6894__A2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5381_ _0787_ _0788_ _0789_ _0523_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7120_ as2650.stack\[4\]\[13\] _2391_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8096__A1 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7843__A1 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7051_ _1518_ _1520_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5004__I _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7071__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7953_ _3191_ as2650.holding_reg\[4\] _3186_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4843__I _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _1099_ _2045_ _2099_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7884_ _3128_ _3111_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7359__C _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8020__B2 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6835_ _0949_ _2044_ _2148_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5909__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8571__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6582__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ _2079_ _2028_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5385__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8505_ _4418_ _3722_ _4335_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5717_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6697_ _1873_ _2012_ _2013_ _1982_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8050__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8436_ _2380_ _3463_ _4429_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5648_ _0982_ _0983_ _1053_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8367_ _2370_ _3589_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ as2650.holding_reg\[4\] _0917_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7318_ _2534_ _2535_ _2559_ _2577_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8087__A1 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8298_ _2712_ _3523_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7834__A1 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6637__A2 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__B _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _1649_ _1278_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5860__A3 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8314__A2 _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5128__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6325__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__A3 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A1 _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4928__I _4433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__I _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A1 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput8 io_in[6] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__7053__A2 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8250__A1 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _4296_ _4345_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4811__A1 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4881_ as2650.cycle\[11\] _0295_ _0311_ _4247_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8553__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6620_ _1920_ _1935_ _1936_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6564__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] _4061_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5502_ _0845_ _0820_ _0742_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5119__A2 as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _1433_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6316__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8221_ _1500_ _4111_ _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5433_ _4137_ _4142_ _4395_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8069__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8152_ _3381_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5364_ _4391_ _0771_ _0772_ _0631_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7103_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7816__A1 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4838__I _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7816__B2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8083_ _1687_ _3314_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _2272_ _2316_ _2327_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A2 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8985_ _0096_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5055__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8792__A2 _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7936_ _3174_ _2365_ _3177_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7867_ _3106_ _3107_ _3108_ _3113_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_54_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8544__A2 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6818_ _2131_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7798_ _3045_ _3006_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6749_ _2007_ _2033_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6307__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6307__B2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8419_ _3555_ _3639_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7807__A1 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__I _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8232__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8783__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6794__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8535__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8299__A1 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8299__B2 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8838__A3 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5263__B _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4658__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8471__A1 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5080_ _0471_ _0499_ _0433_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8574__B _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7969__I as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8223__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7026__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__B2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8990__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5982_ as2650.stack\[1\]\[5\] _1361_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8770_ _2289_ _3925_ _3930_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7721_ as2650.addr_buff\[0\] _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4933_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4864_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7652_ _2685_ _2902_ _2904_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6603_ _1918_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7583_ _2833_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _4302_ _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_59_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7209__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6534_ _0638_ _1849_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6465_ _1781_ _1786_ _1788_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5416_ _0721_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8204_ _3427_ _3428_ _3431_ _1046_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_9184_ _0281_ clknet_leaf_82_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6396_ _1732_ _1733_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8135_ _3319_ _3321_ _3364_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5347_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8066_ _3032_ _3297_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8462__B2 _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ _0367_ _0302_ _0519_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__B _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7017_ as2650.r123_2\[1\]\[3\] _2306_ _2314_ _2310_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6783__I _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8214__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5399__I _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8968_ _0079_ clknet_leaf_15_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7919_ _1259_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8899_ _4041_ _4042_ _3648_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5862__I _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5503__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6551__I1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7256__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8453__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5019__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8756__A2 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6767__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8841__C _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput11 io_in[9] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4580_ _4119_ _4121_ _4123_ _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_122_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6250_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8692__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6298__A3 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _0609_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6181_ _1532_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7247__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5132_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8444__A1 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _0480_ _0481_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6108__I _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8822_ _0424_ _3968_ _3973_ _3974_ _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5012__I _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6758__A1 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8753_ _3901_ _2236_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5965_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5430__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7704_ _2587_ _2955_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__C _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4916_ _0336_ _0340_ _0342_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8684_ _1243_ _3380_ _1782_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5896_ _1272_ _1294_ _1295_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7635_ _0394_ _2884_ _2887_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4847_ _4439_ _4440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7566_ _2554_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4778_ _4093_ _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6930__A1 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6517_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__I _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ _2744_ _2752_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9236_ net47 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8683__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6448_ _1404_ _1771_ _1776_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5497__A1 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6379_ _1716_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9167_ _0264_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8435__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8118_ as2650.stack\[1\]\[2\] _3252_ _3245_ as2650.stack\[0\]\[2\] _1046_ _3349_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8435__B2 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9098_ _0195_ clknet_leaf_82_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8049_ _3168_ _4222_ _4237_ _0388_ _2330_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_102_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8450__A4 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8199__B1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8738__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7410__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__I _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7174__A1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6921__B2 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6688__I _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7477__A2 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9191__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7468__B _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9239__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4701_ _4277_ _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5681_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7165__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7165__B2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8901__A2 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7420_ _2677_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4632_ _4169_ _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6373__C1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6598__I _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _0675_ _0659_ _2608_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4563_ as2650.alu_op\[0\] _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8114__B1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6302_ _0446_ _1495_ _1638_ _1640_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7468__A2 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7282_ _2384_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4494_ as2650.psl\[4\] _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5479__A1 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9021_ _0132_ clknet_leaf_5_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6233_ as2650.stack\[3\]\[8\] _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5007__I _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8417__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6164_ _0383_ _4348_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4846__I _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5115_ _0524_ as2650.cycle\[0\] _0492_ _4245_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ as2650.r123_2\[3\]\[4\] _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6979__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5046_ _4242_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7640__A2 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8805_ _1643_ _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _1330_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_74_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4581__I _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8736_ _0468_ _3884_ _3907_ _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5948_ as2650.stack\[2\]\[3\] _1335_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4757__A3 _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7156__A1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8667_ _2279_ _3859_ _3861_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8353__B1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5879_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7618_ _0441_ _2866_ _2871_ _2714_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5706__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6903__A1 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__C1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8598_ _2762_ _1138_ _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9064__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7549_ _2746_ _2748_ _2747_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8656__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7560__C _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8408__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4693__A2 _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7132__I _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6198__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4491__I as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7147__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8895__A1 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7942__I0 _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4920__A3 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A2 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7042__I _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7622__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _2229_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6851_ _1186_ _1915_ _2134_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5802_ _0625_ _1199_ _1193_ _1005_ _0856_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _1833_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8521_ _3697_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5733_ _4104_ _0959_ _1134_ _1032_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8886__A1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8452_ _1422_ _3660_ _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5664_ _1056_ _1061_ _1063_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7403_ _2630_ _0412_ _2546_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4615_ _4208_ _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8383_ _2903_ _3056_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5595_ _0996_ _0999_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7334_ _2592_ _2538_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4546_ as2650.r123\[1\]\[2\] as2650.r123\[0\]\[2\] as2650.r123_2\[1\]\[2\] as2650.r123_2\[0\]\[2\]
+ _4058_ _4109_ _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_116_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7265_ _2524_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4477_ _4070_ _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5960__I _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8924__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8476__C _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9004_ _0115_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6216_ _1554_ _1563_ _1564_ _1549_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7861__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7196_ as2650.stack\[2\]\[10\] _2462_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7613__A2 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _1437_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8810__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5624__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__B2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _0448_ _4317_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_57 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_79 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7377__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5927__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8719_ _3895_ _3896_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8877__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A3 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8892__A4 _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8629__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5870__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5863__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__A2 as2650.cycle\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8801__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7368__A1 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7368__B2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8565__B1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8565__C2 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6206__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8868__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8947__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7037__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ _4218_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _0353_ _4341_ _0562_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_114_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7843__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5854__A1 _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5606__A1 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _3189_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6903_ _1668_ _2048_ _1818_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7883_ _0310_ _2494_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7359__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6834_ _0950_ _2100_ _1836_ _2147_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8020__A2 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7656__B _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _1989_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6582__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A3 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8504_ _1493_ _0641_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5716_ _4100_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8859__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6696_ _1942_ _1981_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8435_ _2380_ _0463_ _3654_ _0399_ _4424_ _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5647_ _0579_ _1039_ _1052_ _0745_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8366_ _2972_ _2366_ _4435_ _3540_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _4175_ _4396_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8487__B _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7317_ _2563_ _2567_ _2576_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__I _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4529_ _4068_ _4122_ _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8297_ _0392_ _2723_ _3234_ _3522_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9102__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7248_ _4308_ _1481_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5845__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7179_ _2450_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__A4 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__A1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4584__A1 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7522__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5128__A3 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7589__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput9 io_in[7] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4944__I _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8250__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5064__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4811__A2 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4880_ _0309_ _4255_ _4313_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7476__B _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7761__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ _1863_ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5708__C _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5501_ _0817_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7513__A1 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _1798_ _1787_ _1799_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6316__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8220_ _3446_ _3399_ _3447_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5432_ _0585_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9125__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _0764_ _0756_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8151_ as2650.stack\[5\]\[3\] _2455_ _3347_ as2650.stack\[6\]\[3\] _3381_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_114_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7102_ _0706_ _0702_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8082_ _3273_ _3275_ _3312_ _3313_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5294_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ as2650.r123_2\[1\]\[7\] _2304_ _2326_ _2321_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__I _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8326__I _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8241__A2 _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7044__A3 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8984_ _0095_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5055__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _1540_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7866_ _3109_ _2496_ _3110_ _3112_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_35_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6004__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _4098_ _1861_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7797_ _3045_ _3003_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5685__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6748_ _2010_ _2032_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6679_ _1963_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8418_ _3512_ _3627_ _3634_ _3277_ _3238_ _3638_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8349_ _2970_ _3572_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7405__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5818__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__I _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8232__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__I _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6243__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6794__A2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7991__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7743__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7743__B2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9148__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8299__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8471__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5285__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4674__I as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8223__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6234__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5981_ _1309_ _1360_ _1362_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8590__B _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7982__A1 _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7720_ _2970_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4932_ _4346_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7918__C _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7651_ _2903_ _2685_ _2571_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4863_ _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7734__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ _1894_ _1904_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7582_ _2834_ _2835_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ _4387_ _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _1819_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ as2650.stack\[6\]\[8\] _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8203_ as2650.stack\[7\]\[5\] _3246_ _3244_ as2650.stack\[4\]\[5\] _3430_ _3431_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__4849__I _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5415_ _0703_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9183_ _0280_ clknet_leaf_41_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7225__I _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _1690_ _0410_ _1730_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8134_ _0881_ _4135_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5346_ as2650.holding_reg\[1\] _0585_ _0751_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8065_ _3288_ _3296_ _0814_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8462__A2 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5277_ _0674_ _0522_ _0686_ _0668_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7016_ _1932_ _1933_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6285__B _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8214__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8967_ _0078_ clknet_leaf_15_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7918_ _3156_ _3159_ _3160_ _3161_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8898_ _3191_ _4039_ _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ _3079_ _3086_ _3096_ _0306_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A1 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7844__B _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__I as2650.cycle\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A1 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6974__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A2 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__A2 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4494__I as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6767__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__B _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8508__A3 _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7716__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__A1 _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8141__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4669__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8692__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ as2650.carry _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _0782_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7247__A3 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8444__A2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6455__A1 as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5721__C _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _4386_ _4382_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8821_ _1477_ _3968_ _3310_ _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6758__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6833__B _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8752_ _1108_ _3911_ _3912_ as2650.r123\[2\]\[5\] _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ as2650.psu\[2\] _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7703_ _2953_ _2954_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5430__A2 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__B _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ _0336_ _0309_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8683_ _2299_ _3865_ _3870_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5895_ as2650.stack\[3\]\[2\] _1285_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6124__I _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7634_ _2885_ _0412_ _2886_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4846_ _4438_ _4439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__A1 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _2809_ _2819_ _2715_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _4315_ _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4941__A1 _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _1825_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7496_ _2376_ _2745_ _2749_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8132__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9235_ net47 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4579__I _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ as2650.stack\[0\]\[10\] _1774_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6694__A1 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5497__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9166_ _0263_ clknet_leaf_4_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6378_ _0881_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8495__B _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8117_ as2650.stack\[3\]\[2\] _2388_ _3347_ as2650.stack\[2\]\[2\] _3348_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_142_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8435__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5329_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9097_ _0194_ clknet_leaf_82_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8048_ _2582_ _3279_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5631__C _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8199__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7558__C _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5421__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5359__B _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__I _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8371__A1 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__I _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8980__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7229__A3 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__I0 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _4293_ _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5680_ _1055_ _1010_ _1081_ _0941_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__8362__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ _4223_ _4224_ _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5783__I _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6373__B1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__C2 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7350_ _0676_ _0659_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4562_ _4155_ _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _4371_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7281_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4493_ _4082_ _4084_ _4086_ _4059_ _4087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9020_ _0131_ clknet_leaf_74_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6232_ _1576_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8417__A2 _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6163_ _1509_ _4317_ _1511_ _1516_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5114_ _4064_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _1453_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6119__I _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _0432_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7659__B _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7928__A1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8804_ _3939_ _3940_ _3957_ _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6996_ _2297_ _2292_ _2298_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8735_ _1466_ _0570_ _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5947_ _1294_ _1334_ _1338_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8666_ as2650.stack\[6\]\[0\] _3860_ _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8353__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ _4364_ _0479_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8353__B2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7617_ _2587_ _2869_ _2870_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6364__B1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4829_ _4270_ _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6364__C2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8597_ _3808_ _3809_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7548_ _1020_ _1015_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8105__A1 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7479_ _1304_ net11 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8656__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6667__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9149_ _0246_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8509__I _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__I _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6192__C _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8592__A1 _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8344__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7147__A2 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5158__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8895__A2 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7942__I1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8847__C _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5330__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7323__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5633__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__B _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8032__B1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _2161_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _1201_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__A1 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6781_ _1850_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8520_ _2410_ _3308_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5732_ _0799_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5149__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8451_ as2650.pc\[14\] _3669_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5663_ _1066_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7402_ _2634_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6897__A1 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _4146_ _4152_ _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8382_ _3603_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ _0996_ _0999_ _0930_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7333_ net30 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4545_ _4138_ _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8638__A2 _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5018__I _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__A1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7264_ _2523_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4476_ _4066_ as2650.ins_reg\[1\] _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7310__A2 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9003_ _0114_ clknet_leaf_44_wb_clk_i as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6215_ net20 _1559_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4857__I _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5321__A1 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _2459_ _1396_ _2463_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6146_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _1437_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8810__A2 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8492__C _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5624__A2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input10_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__I _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__B1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_58 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9100__D _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7377__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8574__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ _2285_ _2282_ _2286_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8718_ _3892_ _2312_ _3893_ _0901_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8649_ _1781_ _3848_ _3850_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8877__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__I _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6888__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9181__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A4 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4767__I _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5863__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8262__B1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7299__B _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5598__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8014__B1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8565__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8565__B2 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8317__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8868__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6879__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5551__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8149__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ as2650.pc\[8\] _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7988__I _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7056__A1 _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7951_ _1018_ _3176_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9054__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7002__B _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6902_ _4204_ _1837_ _2213_ _2047_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7882_ _2352_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5301__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8556__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6833_ _2144_ _2102_ _1818_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ as2650.r0\[3\] _4089_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5385__A4 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8503_ _0566_ _3718_ _3719_ _3720_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_91_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5715_ as2650.r123\[0\]\[6\] _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6695_ _4098_ _1875_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8859__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8434_ _1422_ _0392_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5646_ _0742_ _1050_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_104_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8365_ _0399_ _3585_ _3581_ _2597_ _3587_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5577_ _0577_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7316_ _2541_ _2347_ _2570_ _2573_ _2575_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4528_ as2650.r123\[1\]\[4\] as2650.r123\[0\]\[4\] as2650.r123_2\[1\]\[4\] as2650.r123_2\[0\]\[4\]
+ _4058_ _4110_ _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8296_ _2552_ _3521_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6288__B _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4587__I _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7247_ _2503_ _2504_ _2505_ _2506_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4459_ _4052_ _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7178_ _2446_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7047__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__B1 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _0437_ _4235_ _1477_ _1480_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__C1 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5781__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A2 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5086__C _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7522__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4497__I _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5836__A2 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7589__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8786__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7757__B _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6549__B1 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8914__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5500_ _0902_ _0903_ _0904_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_119_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ as2650.stack\[6\]\[13\] _1785_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7513__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8710__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6316__A3 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5431_ _0636_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6572__I0 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8150_ _3379_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5362_ _0764_ _0756_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _2385_ _2363_ _2386_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8081_ _3268_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5293_ _0700_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7032_ _1961_ _1996_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7511__I _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A4 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8983_ _0094_ clknet_leaf_69_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5055__A3 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6127__I _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ _3175_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8529__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7865_ _0411_ _2712_ _3111_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__A1 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6004__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _2129_ _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7796_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _1998_ _2035_ _2062_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_56_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _1964_ _1994_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5629_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8417_ _0425_ _3636_ _3637_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5515__A1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8348_ _2972_ _2720_ _3540_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7268__A1 _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8279_ as2650.stack\[5\]\[7\] _3242_ _3251_ as2650.stack\[6\]\[7\] _3505_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8517__I _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7421__I _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8768__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7440__A1 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4780__I _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7743__A2 _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5754__A1 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6951__B1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6554__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7259__A1 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5116__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4955__I _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8759__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A1 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7431__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ as2650.stack\[1\]\[4\] _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7982__A2 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4931_ _0355_ _0293_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5993__A1 _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7650_ _2536_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4862_ _4352_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7734__A2 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6601_ _1913_ _1917_ _1912_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7581_ _1093_ _1103_ _2797_ _2756_ _2798_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5745__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4793_ _4386_ _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _0651_ _1834_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _1785_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8111__B _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7506__I _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8202_ _3429_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5414_ as2650.stack\[7\]\[9\] _0821_ _0822_ as2650.stack\[6\]\[9\] _0823_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9182_ _0279_ clknet_leaf_41_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _0477_ _1494_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_115_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8133_ _3361_ _3362_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0753_ _0539_ _4394_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8064_ _0360_ _3291_ _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _0676_ _0682_ _0684_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7015_ _2111_ _2302_ _2313_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_68_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__C _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8214__A3 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__A2 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8966_ _0077_ clknet_leaf_43_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7917_ _1507_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8897_ _4023_ _4037_ as2650.psu\[4\] _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ _3069_ _2959_ _3095_ _2861_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4539__A2 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _3009_ _2768_ _2335_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6320__I _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5364__C _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6161__A1 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A2 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6464__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4475__A1 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6216__A2 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7413__A1 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5019__A3 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9115__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7716__A2 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7326__I _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4950__A2 _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8141__A2 _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6230__I _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__C _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5130_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6455__A2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _4378_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7404__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8820_ _1510_ _3972_ _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8751_ _0551_ _0740_ _2198_ _3918_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_52_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5966__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5963_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7702_ _2936_ _2951_ _2952_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4914_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5894_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8682_ as2650.stack\[6\]\[7\] _3866_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7945__B _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7633_ _2545_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _4253_ _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7564_ _2817_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7664__C _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4776_ _4369_ _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _1831_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7495_ _2745_ _2750_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4941__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8132__A2 _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6140__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9234_ net47 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6446_ _1396_ _1771_ _1775_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7891__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9165_ _0262_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6377_ as2650.psl\[1\] _1713_ _1658_ _1660_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8116_ _1572_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5328_ _4398_ _0482_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_103_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9096_ _0193_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__A1 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8047_ _1274_ _4268_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6446__A2 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9138__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8199__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8949_ _0060_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5957__A1 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6315__I _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5709__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8371__A2 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6382__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7229__A4 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8705__I _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A1 _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8362__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4630_ as2650.psl\[6\] _4060_ _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6373__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6373__B2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _4148_ _4154_ _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8114__A2 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6300_ _0677_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7280_ net29 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6125__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4492_ _4085_ _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8596__B _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6231_ _1576_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _4320_ _0364_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_124_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7625__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5113_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ as2650.r123_2\[3\]\[3\] _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5304__I _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__B1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ _0461_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7928__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8803_ _0423_ _1462_ _3942_ _3194_ _3956_ _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_93_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6995_ as2650.stack\[5\]\[6\] _2293_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8734_ _1729_ _1132_ _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5946_ as2650.stack\[2\]\[2\] _1335_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4611__A1 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8665_ _3858_ _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8353__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _2832_ _2715_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4828_ _4421_ _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6364__A1 _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__B2 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8596_ _1312_ _3750_ _2482_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4759_ as2650.cycle\[13\] _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7547_ _1490_ _2745_ _2744_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6116__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7478_ _0335_ _2734_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7864__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ _4341_ _1245_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__C _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9148_ _0245_ clknet_leaf_46_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7616__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__A2 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9079_ _0176_ clknet_leaf_19_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7569__C _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4850__A1 _4440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8592__A2 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4602__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8260__I _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5158__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__A1 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__A2 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4963__I _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4841__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__C _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8032__B2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8583__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5800_ _1164_ _1167_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6780_ _1832_ _2061_ _2095_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5397__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5731_ _1082_ _4102_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5662_ _0994_ _1002_ _0992_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6346__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5149__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8450_ _3650_ _3068_ _1407_ _3602_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7401_ _2588_ _2589_ _2635_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4613_ _4206_ _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8381_ _1407_ _3602_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6897__A2 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5593_ _0924_ _0934_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _2587_ _2590_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8099__A1 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4544_ as2650.r0\[2\] _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7263_ _2496_ _2499_ _2500_ _2522_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__7846__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4475_ _4065_ _4068_ _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9002_ _0113_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6214_ _1312_ _1555_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7194_ as2650.stack\[2\]\[9\] _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5321__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6145_ net1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_112_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__I _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8271__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _1300_ _1438_ _1443_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5969__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5027_ _4277_ _4381_ _4056_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A1 _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8023__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_59 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8574__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8970__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6978_ as2650.stack\[5\]\[1\] _2283_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8717_ as2650.r123\[1\]\[2\] _3890_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8648_ as2650.stack\[7\]\[8\] _3849_ _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8877__A3 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6888__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8579_ _2376_ _1670_ _3791_ _3792_ _0380_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4899__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5863__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__I _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4783__I _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4823__A1 _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8014__B2 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6576__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8868__A3 _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5000__A1 _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7828__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6500__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A3 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8253__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7056__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A1 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6803__A2 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8993__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7950_ _3188_ _2377_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4814__A1 _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6901_ _1094_ _2049_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7002__C _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7881_ _2498_ _3126_ _2342_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_78_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _4212_ _1837_ _2145_ _2047_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6763_ _2024_ _2027_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__B _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8308__A2 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8502_ _4170_ _2343_ _1630_ _1248_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5714_ _1054_ _0983_ _1118_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6694_ _4099_ _1890_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8433_ _2597_ _3652_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5645_ _1018_ _0734_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8364_ _2369_ _3027_ _3586_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5576_ as2650.r123\[0\]\[4\] _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7819__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7315_ _4409_ _2539_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4868__I _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4527_ _4071_ _4120_ _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8295_ _2584_ _4073_ _3520_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8492__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7246_ _4322_ _4329_ _1253_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4458_ as2650.ins_reg\[4\] _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8492__B2 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ _2247_ _2419_ _2437_ _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7047__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8244__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6128_ _4243_ _4445_ _0449_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5699__I _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A1 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ as2650.r123_2\[0\]\[6\] _1376_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__A1 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A2 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__B1 _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5781__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A3 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8180__B1 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5533__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6730__A1 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7090__S _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8786__A2 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8713__I _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6549__B2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8588__C _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8710__A2 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _4191_ _4377_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6572__I1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _0628_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7100_ _4432_ _2359_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8080_ _3299_ _3301_ _3311_ _3273_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_142_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7999__I _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9021__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7031_ _2247_ _2316_ _2325_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__A1 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8982_ _0093_ clknet_3_1__leaf_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5312__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6788__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9171__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout53_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7933_ _2407_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5460__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7864_ _1481_ _0552_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _1968_ _1858_ _4090_ as2650.r0\[4\] _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7795_ as2650.addr_buff\[3\] _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7752__A3 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _2002_ _2034_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6677_ _1966_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8701__A2 _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8416_ _0425_ _3626_ _1622_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5628_ _1032_ _1012_ _1013_ _0871_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4598__I _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8347_ _3238_ _3570_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9106__D _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5559_ _0808_ _0948_ _0965_ _0694_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7268__A2 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8465__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8278_ as2650.stack\[1\]\[7\] _2456_ _3380_ as2650.stack\[0\]\[7\] _1047_ _3504_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_104_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _0465_ _2485_ _2487_ _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_105_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__B2 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6951__B2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8153__B1 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4502__S _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6703__A1 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__I1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7259__A2 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8456__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8208__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8759__A2 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__I _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5442__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4971__I _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4861_ _4446_ _0291_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7195__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7059__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6600_ _1914_ _1916_ _1899_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_53_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7580_ _1093_ _1103_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5745__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ _4239_ _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4953__B1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6531_ _0659_ _1835_ _1833_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6462_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8111__C _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8201_ as2650.stack\[5\]\[5\] _3241_ _1572_ as2650.stack\[6\]\[5\] _3429_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5413_ _0717_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6393_ _1707_ _1721_ _1728_ _1730_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_9181_ _0278_ clknet_leaf_45_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8132_ _0952_ _4130_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5344_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_82_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8063_ _0787_ _3292_ _3293_ _2366_ _3294_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _0521_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7014_ as2650.r123_2\[1\]\[2\] _2306_ _2312_ _2310_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__I _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8214__A4 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8965_ _0076_ clknet_leaf_63_wb_clk_i as2650.r123_2\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A1 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7916_ _0596_ _3156_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_37_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7397__C _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8896_ _4038_ _4040_ _3648_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7847_ _2886_ _3090_ _3094_ _4406_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7778_ _2555_ _2370_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6933__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _1817_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6161__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4711__A3 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7110__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__A4 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8610__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5887__I _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7607__I _4440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8677__A1 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8429__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4966__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7101__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__I _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _4372_ _0472_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8882__B _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7404__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8601__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6612__B1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8750_ _1039_ _3911_ _3909_ as2650.r123\[2\]\[4\] _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _0708_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7701_ _2951_ _2952_ _2936_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ as2650.cycle\[8\] _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8681_ _2297_ _3865_ _3869_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8365__B1 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5893_ _0845_ _1292_ _1281_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7632_ net54 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4844_ _4436_ _4437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__B _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7563_ _2735_ _2775_ _2791_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _4293_ _4324_ _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8117__B1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6514_ _1830_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8668__A1 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7494_ _2746_ _2748_ _2747_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__A3 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ as2650.stack\[0\]\[9\] _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7340__A1 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8927__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6143__A2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9164_ _0261_ clknet_leaf_79_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7891__A2 _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6376_ _0549_ _1021_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8115_ as2650.stack\[5\]\[2\] _3252_ _3245_ as2650.stack\[4\]\[2\] _0905_ _3346_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5327_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9095_ _0192_ clknet_3_0__leaf_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8046_ _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8792__B _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5654__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8948_ _0059_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7159__A1 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8879_ _1622_ _1495_ _4026_ _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7159__B2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6331__I _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__B _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7634__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5645__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6070__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4471__I2 as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8898__A1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7337__I _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _4153_ _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5285__C _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4491_ as2650.ins_reg\[1\] _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6125__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6676__A3 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4687__A2 as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4696__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ _4241_ _1512_ _1248_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_97_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5112_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _1452_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8822__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7800__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7389__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8802_ _3133_ _3946_ _3950_ _3955_ _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5939__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _1324_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6061__A1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8733_ _1238_ _3883_ _3905_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5945_ _1290_ _1334_ _1337_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4611__A2 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8889__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8664_ _3858_ _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5876_ _4045_ _1247_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_139_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7615_ _2854_ _2868_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _4417_ _4418_ _4420_ _4351_ _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8595_ _3798_ _3807_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6364__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7546_ _2562_ _2800_ _0326_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4758_ _4340_ _4351_ _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7477_ net55 _2581_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7313__A1 _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4689_ as2650.cycle\[4\] _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_88_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6428_ _1762_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7864__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9147_ _0244_ clknet_leaf_34_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__A2 _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8813__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9078_ _0175_ clknet_leaf_22_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8029_ _0414_ _3259_ _3261_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7585__C _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5386__B _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6107__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7855__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5866__A1 _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5405__I _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8804__A1 _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6815__B1 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6291__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__A2 _4433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__A1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7791__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6594__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _4185_ _1079_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5661_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7067__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5149__A3 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _2347_ _2632_ _2638_ _2657_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4612_ _4205_ _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9128__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8380_ _1399_ _3580_ _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5554__B1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5592_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7331_ _2588_ _2589_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8099__A2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _4136_ _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5306__B1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7262_ _2480_ _2507_ _2508_ _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_132_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7846__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4474_ _4067_ _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5306__C2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9001_ _0112_ clknet_leaf_46_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6213_ _1561_ _1556_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7193_ _2457_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _1488_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8271__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ as2650.stack\[0\]\[3\] _1439_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6282__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6282__B2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5026_ _4313_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6409__I0 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8559__B1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6146__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4832__A2 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8023__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _1289_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8716_ _3891_ _3894_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4596__A1 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _1319_ _1273_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8647_ _3847_ _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5859_ _4439_ _0341_ _0442_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8877__A4 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8578_ _1550_ _1650_ _0793_ _1561_ _1670_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_120_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7529_ _2740_ _2581_ _1687_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A1 _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7065__A3 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8262__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__A2 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8014__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__A1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6500__A2 _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A4 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4974__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8253__A2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5067__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8890__B _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A2 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _1104_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7880_ _4048_ _4415_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6016__A1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _0953_ _1813_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6567__A2 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6762_ _2076_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8308__A3 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8501_ _3168_ _1643_ _0553_ _1635_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5713_ _0579_ _1108_ _1117_ _0745_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7516__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6693_ _1976_ _2008_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8432_ _3650_ _3651_ _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5644_ _0817_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8363_ _2370_ _2355_ _4428_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5575_ _0912_ _0578_ _0981_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7525__I _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7314_ _4048_ _1509_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4750__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4526_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _4109_ _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8294_ _2898_ _4096_ _3469_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7245_ _4441_ _1481_ _1459_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5045__I _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ _4050_ _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8492__A2 _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _2321_ _2422_ _2423_ _1319_ _2447_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6127_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__A2 _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6058_ _1429_ _1382_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__A2 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5009_ _0428_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6007__A1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4584__A4 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6540__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8180__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8180__B2 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6730__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4794__I _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7746__A1 _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8215__B _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6549__A2 _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6514__I _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5221__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8171__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4969__I _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6389__C _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4732__A1 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5360_ _0767_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8885__B _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5291_ as2650.psu\[1\] _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8474__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6485__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7030_ as2650.r123_2\[1\]\[6\] _2304_ _2324_ _2321_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7080__I _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8981_ _0092_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6788__A2 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7932_ _2473_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _4416_ _0315_ _2495_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7737__A1 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _2083_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7794_ _3040_ _3042_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5212__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6745_ _2058_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6960__A2 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7683__C _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _1976_ _1980_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8162__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8415_ _3068_ _2537_ _3635_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5627_ _0951_ _0872_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8346_ _3441_ _3563_ _3564_ _3569_ _1488_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4723__A1 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _0692_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _4102_ _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8465__A2 _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8277_ as2650.stack\[3\]\[7\] _2389_ _1574_ as2650.stack\[2\]\[7\] _3503_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5489_ _0528_ _0543_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _4353_ _1477_ _0291_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8217__A2 _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7159_ _2421_ _2422_ _2423_ _0969_ _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_59_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9122__D _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6779__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7728__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6334__I _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5203__A2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6400__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6951__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4789__I _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7900__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6703__A2 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_7_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_69_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__I _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__I _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6219__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7416__B1 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5993__A3 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _4331_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _4328_ _4384_ _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ _1806_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4953__A1 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4953__B2 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4699__I _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8695__A2 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8200_ as2650.stack\[1\]\[5\] _2455_ _3379_ as2650.stack\[0\]\[5\] _0721_ _3428_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_5412_ _0713_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9180_ _0277_ clknet_3_2__leaf_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6392_ _1729_ _1469_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8131_ _0952_ _4130_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5343_ _4150_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8062_ _0375_ _3274_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5274_ _4216_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7013_ _1928_ _1930_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5323__I _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8634__I _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8964_ _0075_ clknet_leaf_61_wb_clk_i as2650.r123_2\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6630__A1 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5433__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7915_ _2382_ _2478_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8895_ _3197_ _4039_ _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7846_ _3069_ _2531_ _3093_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8383__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7694__B _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7777_ _2863_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _1821_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _1967_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__9117__D _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6697__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6161__A3 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8329_ _2385_ _2955_ _3553_ _1489_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5121__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6329__I _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9011__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8126__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5408__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8429__A2 _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7101__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4546__S0 _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6860__A1 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7779__B _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4982__I _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8601__A2 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6612__B2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _1269_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7700_ _2735_ _2775_ _2790_ _2937_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_4912_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8680_ as2650.stack\[6\]\[6\] _3866_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5892_ as2650.pc\[2\] _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8365__A1 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8365__B2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7631_ _2881_ _2883_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4843_ _4435_ _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7562_ _2788_ _1091_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4926__A1 _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ _4367_ _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8117__B2 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8122__C _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _1729_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7493_ _2746_ _2747_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _1769_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9163_ _0260_ clknet_leaf_77_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6375_ _1712_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7891__A3 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8114_ as2650.stack\[7\]\[2\] _3250_ _3251_ as2650.stack\[6\]\[2\] _3345_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ _4357_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9094_ _0191_ clknet_leaf_82_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8045_ _4423_ _3276_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__S0 _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5257_ _0666_ _4307_ _0519_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5053__I _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__A2 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5188_ _0596_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5988__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4892__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8947_ _0058_ clknet_leaf_50_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9034__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8356__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8878_ _0480_ _3208_ _4025_ _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7829_ net53 _3076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6906__A2 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5656__C _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9184__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8659__A2 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5342__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8539__I _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__S0 _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8831__A2 _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5898__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8595__A1 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8347__A1 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8898__A2 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__B1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ as2650.r123\[1\]\[6\] _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7353__I _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _4345_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8893__B net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7086__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _4438_ _0519_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4519__S0 _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ as2650.r123_2\[3\]\[2\] _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8822__A2 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ as2650.cycle\[13\] _4447_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9057__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8586__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8801_ _1630_ _3954_ _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _2295_ _2292_ _2296_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8732_ _3885_ _2326_ _3888_ as2650.r123\[1\]\[7\] _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5944_ as2650.stack\[2\]\[1\] _1335_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8663_ _1436_ _1349_ _2280_ _1347_ _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_90_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5875_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7614_ _2867_ _2817_ _2857_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4826_ _4381_ _4303_ _4419_ _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8594_ _4204_ _0466_ _3806_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7972__B net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7545_ _1501_ _1104_ _2799_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4757_ _4342_ _4343_ _4350_ _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5048__I _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7476_ _2709_ _2732_ _2675_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ as2650.cycle\[5\] _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8510__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8359__I _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _1678_ _1751_ _1759_ _0437_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5324__A1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9146_ _0243_ clknet_leaf_34_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6358_ _4450_ _4306_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7077__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5309_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9077_ _0174_ clknet_leaf_19_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _1524_ _1626_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_88_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6824__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8028_ _3222_ _3260_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5511__I _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_21_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_leaf_21_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6543__S _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8329__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8501__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__I _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8265__B1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8804__A2 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__B2 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__I _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7240__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8917__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6043__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7791__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _1062_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8888__B as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7543__A2 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4611_ _4129_ _4132_ _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5554__A1 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ as2650.holding_reg\[3\] _4378_ _0915_ _0921_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_129_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7330_ as2650.pc\[1\] net8 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4542_ _4071_ _4135_ _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7261_ _2511_ _2514_ _2517_ _2520_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_128_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7083__I _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _4066_ as2650.ins_reg\[1\] _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_89_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9000_ _0111_ clknet_leaf_53_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6212_ _1055_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _2459_ _1386_ _2461_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _1492_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _1294_ _1438_ _1442_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6282__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _4325_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8559__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8559__B2 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6409__I1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4832__A3 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6976_ _2279_ _2282_ _2284_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8715_ _3892_ _2309_ _3893_ _0811_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4596__A2 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ _1322_ _1280_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _0337_ _4245_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8646_ _3847_ _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8731__A1 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4809_ _4371_ _4385_ _4399_ _4402_ _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5789_ _1191_ _1184_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8577_ _3787_ _3788_ _3789_ _3790_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_135_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7528_ _2707_ _2765_ _2783_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7459_ _2634_ _2659_ _2704_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5506__I _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A2 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9129_ _0226_ clknet_leaf_33_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8798__A1 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6273__A2 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6337__I _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5241__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7222__A1 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6025__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8722__A1 as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6328__A3 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8501__B _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7289__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9035__D _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6956__B _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8789__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7461__A1 _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4814__A3 _4407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7213__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _0951_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _2023_ _2030_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7078__I _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5712_ _0742_ _1115_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8500_ _2352_ _1512_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6692_ _1980_ _1992_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7516__A2 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5643_ _0831_ _1042_ _1045_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8431_ _3068_ _1407_ _3602_ _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8362_ _1693_ _3024_ _3584_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5754__C _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5574_ _0571_ _0968_ _0971_ _0980_ _0576_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7313_ _4336_ _2571_ _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4525_ _4118_ _4078_ _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8293_ _3441_ _3514_ _3518_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4750__A2 as2650.cycle\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5326__I _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _0353_ _4346_ _0556_ _1513_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _4049_ _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8229__B1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7175_ _1128_ _2409_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_63_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _0550_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6255__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6057_ as2650.pc\[14\] _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__I _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__A3 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ _4296_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6959_ _2043_ _2268_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8629_ _2285_ _3834_ _3837_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8180__A2 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6067__I _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5855__B _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6557__I0 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7626__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8171__A2 _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5574__C _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4732__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__I _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5290_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7682__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6485__A2 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7361__I _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7434__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8980_ _0091_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7931_ _0584_ _3166_ _3173_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7862_ _2512_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7737__A2 _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ as2650.r0\[5\] _4089_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _3015_ _3019_ _3041_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _0775_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6675_ _1983_ _1991_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8162__A2 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__I _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8414_ _2384_ _3088_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5626_ _0655_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6173__A1 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8345_ _3475_ _3566_ _3561_ _2595_ _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5557_ _0958_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5056__I _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4508_ _4095_ _4097_ _4101_ _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8276_ _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _0893_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7673__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__I _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7227_ _4323_ _1253_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _0978_ _2428_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _1463_ _0369_ _1264_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7089_ as2650.addr_buff\[4\] _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__B _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8153__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7900__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7664__A1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7664__B2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7416__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7416__B2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9090__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7784__C _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _4298_ _4380_ _4383_ _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_82_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4953__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8144__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6460_ _1346_ _1782_ _1783_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8896__B _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _0816_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6391_ _4248_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8130_ _2710_ _3359_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5342_ _4147_ _4153_ _0598_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8061_ _4345_ _4434_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7655__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ _0681_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7012_ _2061_ _2302_ _2311_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7407__A1 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8963_ _0074_ clknet_3_5__leaf_wb_clk_i as2650.r123_2\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7914_ _3156_ _3157_ _3158_ _2629_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_3_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__A1 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8894_ _4051_ _1497_ _4037_ _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7845_ _4436_ _3077_ _3091_ _3092_ _2989_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_54_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8650__I _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5197__A2 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7776_ _1694_ _3024_ _3025_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4988_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6727_ _1806_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6170__I _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6658_ _1971_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7894__A1 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5609_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_46_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6589_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6161__A4 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8328_ _1380_ _2538_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7646__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8259_ _3472_ _3482_ _3485_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5121__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4880__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6621__A2 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A2 _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8950__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A3 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8126__A2 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6137__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7885__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7637__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4546__S1 _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8062__A1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6612__A2 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _0700_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5891_ _1272_ _1290_ _1291_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8365__A2 _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8470__I _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7630_ _2854_ _2868_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4842_ _4434_ _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7561_ _2528_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4773_ _4294_ _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4926__A2 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8117__A2 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6128__A1 _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6512_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7492_ _1019_ _1014_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_134_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6443_ _1386_ _1771_ _1773_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6374_ _0784_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_9162_ _0259_ clknet_leaf_71_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5325_ _0698_ _0730_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8113_ _3343_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9093_ _0190_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5639__B1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5256_ _0630_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8044_ _4221_ _4237_ _0812_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4537__S1 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6851__A2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8645__I _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ as2650.idx_ctrl\[0\] _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4862__A1 _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8973__CLK clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8946_ _0057_ clknet_leaf_59_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A1 _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8877_ _0432_ _1509_ _2498_ _2989_ _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_7828_ net40 _3051_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6367__A1 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ net39 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4917__A2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5342__A2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7619__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8292__A1 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8292__B2 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__S1 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__I _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__A1 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8044__A1 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A1 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A1 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5030__A1 _4437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__B2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7858__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _0370_ _4305_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8283__A1 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7086__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _1451_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4519__S1 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5041_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8996__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8586__A2 _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8800_ _3700_ _3951_ _3953_ _4308_ _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6597__A1 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6992_ as2650.stack\[5\]\[5\] _2293_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8731_ _1179_ _3883_ _3904_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5943_ _1284_ _1334_ _1336_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8662_ _1800_ _3849_ _3857_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6349__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5874_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _2735_ _2775_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _4249_ _4419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _1490_ _3754_ _0365_ _1028_ _3805_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5329__I _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7544_ _2797_ _2756_ _2798_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7972__C _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4756_ _4290_ _4346_ _4349_ _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_105_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5572__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7849__A1 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7849__B2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7475_ _2710_ _2529_ _2730_ _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4687_ _4264_ as2650.cycle\[11\] _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8510__A2 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6426_ _0476_ _1759_ _1760_ _1761_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9145_ _0242_ clknet_leaf_30_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _1639_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7077__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9076_ _0173_ clknet_leaf_19_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _4320_ _4399_ _0564_ _1478_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_130_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9001__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8027_ _2471_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _0646_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_112_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8026__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8929_ _0040_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8329__A2 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_3_5__leaf_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__I1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7454__I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8501__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5079__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__B _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A1 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__C _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7240__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6533__I _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7565__S _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _4201_ _4202_ _4203_ _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5590_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6751__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4988__I _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4541_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _4109_ _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7260_ _4276_ _2332_ _2519_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4472_ as2650.ins_reg\[0\] _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5306__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6503__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6211_ _1554_ _1558_ _1560_ _1549_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9024__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7191_ as2650.stack\[2\]\[8\] _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8256__A1 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ as2650.stack\[0\]\[2\] _1439_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__I _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9174__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5024_ _0438_ _0442_ _0443_ _4266_ _4275_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8559__A2 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8144__B _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ as2650.stack\[5\]\[0\] _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8714_ _3886_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5926_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6990__A1 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8645_ _3846_ _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5857_ _0527_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8731__A2 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4808_ _4401_ _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8576_ _1865_ _0502_ _1701_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6742__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5788_ _1189_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7527_ _1305_ _2583_ _2780_ _2782_ _2675_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _4263_ as2650.cycle\[1\] _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7274__I _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__A2 _4437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8495__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7458_ _2585_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6409_ _1690_ _1746_ _1648_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7389_ _2639_ _2614_ _2646_ _2571_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8247__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9128_ _0225_ clknet_leaf_34_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8798__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9059_ _0156_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__S _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7222__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6353__I _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8183__B1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8722__A2 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8501__C _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9047__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8238__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8789__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7997__B1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7461__A2 _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8410__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5224__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5224__B2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ _2026_ _2029_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6972__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8899__B _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _1088_ _0734_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6691_ _1980_ _1992_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8430_ as2650.pc\[13\] _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5642_ as2650.stack\[5\]\[12\] _0824_ _0827_ as2650.stack\[4\]\[12\] _1047_ _1048_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__8411__C _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8361_ _3000_ _0411_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5573_ _0743_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4511__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7312_ _2568_ _0651_ _2328_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4524_ _4117_ _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8292_ _3475_ _3510_ _3517_ _4048_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7243_ _0739_ _1279_ _2338_ _2502_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4455_ _4048_ _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8229__A1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8229__B2 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5770__C _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7174_ as2650.r123_2\[0\]\[6\] _2420_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _1479_ _0855_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6255__A3 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _1387_ _1427_ _1428_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5007_ _4294_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4805__A4 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8401__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7204__A2 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6958_ _1210_ _2044_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _1305_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6889_ _4202_ _2048_ _2100_ _2201_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8628_ as2650.stack\[7\]\[1\] _3835_ _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6715__A1 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8321__C _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8559_ _1915_ _1472_ _3386_ _0489_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7140__A1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6348__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__I _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7400__C _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5206__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6954__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5509__A2 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6557__I1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8459__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4732__A3 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7682__A2 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7434__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8631__A1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7930_ _3166_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _2489_ _2499_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4506__I _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6812_ _2125_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7792_ _2999_ _1142_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6945__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _0565_ _1812_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8422__B _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6721__I _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8698__A1 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6674_ _1987_ _1990_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _1416_ _3633_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5625_ _1018_ _0779_ _1030_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7980__C _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8344_ _3287_ _3567_ _0357_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5556_ _0780_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ _4100_ _4079_ _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8275_ _1327_ _3500_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5487_ _4144_ _0649_ _0894_ _0646_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_7226_ _4353_ _2486_ _1629_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7673__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8870__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ _2432_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5072__I _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6108_ _0814_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8622__A1 _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7088_ _2376_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6039_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8689__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6164__A2 _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7900__A3 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7113__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8861__A1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6078__I _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7416__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__B _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__I _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4953__A3 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7352__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _0753_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6390_ _4388_ _0621_ _1722_ _1727_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5341_ _4208_ _0602_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8468__I _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7372__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8301__B1 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7655__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8060_ _0462_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8852__A1 _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5272_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5666__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7011_ as2650.r123_2\[1\]\[1\] _2306_ _2309_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5666__B2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7407__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8962_ _0073_ clknet_3_5__leaf_wb_clk_i as2650.r123_2\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5620__I _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7913_ _0597_ _3156_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8893_ _3196_ _4037_ net28 _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7844_ net53 _2821_ _2721_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7775_ _3009_ _0393_ _2546_ _0423_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6394__A2 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__C _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _1836_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6657_ _4159_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7343__A1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ _4125_ _1010_ _1012_ _0804_ _1013_ _0892_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__7894__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6588_ _1902_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8327_ _3487_ _0730_ _3551_ _3532_ _3495_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5539_ _4191_ _0869_ _4206_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__I _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6400__B _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__C _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7646__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8258_ _3310_ _3484_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8843__A1 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_wb_clk_i clknet_3_2__leaf_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8189_ _3416_ _3417_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__A2 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6082__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8126__A3 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7334__A1 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6137__A2 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7885__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8062__A2 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5820__A1 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ as2650.stack\[3\]\[1\] _1285_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ _4265_ _4433_ _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7573__A1 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6376__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7573__B2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _0406_ _2794_ _2813_ _2814_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4772_ _4365_ _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6511_ _0549_ _0559_ _1806_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_53_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7491_ _2736_ _2679_ _2641_ _2642_ _2681_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__6128__A2 _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6442_ as2650.stack\[0\]\[8\] _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7876__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_opt_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9161_ _0258_ clknet_leaf_73_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8198__I _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6373_ as2650.psl\[7\] _1214_ _1708_ _0610_ _0609_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_8112_ _4294_ _0445_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _0733_ _0547_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9092_ _0189_ clknet_leaf_81_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8043_ _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5255_ _0663_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5186_ as2650.idx_ctrl\[1\] _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8589__B1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8945_ _0056_ clknet_leaf_59_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4614__A2 _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8876_ _0486_ _1461_ _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7827_ _2686_ _3072_ _3074_ _2929_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7564__A1 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6367__A2 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ _2929_ _3004_ _3007_ _2686_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _1948_ _2024_ _2025_ _1988_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7316__A1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7689_ _2936_ _2939_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8610__B _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7867__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A1 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5342__A3 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7619__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8816__A1 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6557__S _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6356__I _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4853__A2 _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8044__A2 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__B2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7004__B1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7555__A1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6358__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8752__B1 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5030__A2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7307__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7858__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8807__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8283__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ as2650.addr_buff\[7\] _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_111_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8035__A2 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5170__I _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7243__B1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6991_ _1316_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7794__A1 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6597__A2 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8730_ _3885_ _2324_ _3888_ as2650.r123\[1\]\[6\] _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ as2650.stack\[2\]\[0\] _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8661_ as2650.stack\[7\]\[14\] _3847_ _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5873_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7546__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7612_ _2666_ _2850_ _2862_ _2865_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ as2650.cycle\[9\] _4335_ _4338_ _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8592_ _3726_ _3804_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7543_ _1020_ _1034_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4755_ _4348_ _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7474_ _2528_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4686_ _4277_ _4279_ _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7046__B _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6425_ _1754_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9144_ _0241_ clknet_leaf_30_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6356_ _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5307_ _0707_ _0702_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9075_ _0172_ clknet_leaf_19_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6287_ _0546_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6285__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8026_ _1693_ _2539_ _3228_ _3169_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5238_ _0596_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6176__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8026__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5169_ _0571_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8928_ _0039_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7537__A1 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8859_ _3195_ _1476_ _1503_ _3770_ _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5720__B1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8265__A2 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7776__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7528__A1 _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9049__D _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6200__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7645__I _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6751__A2 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _4133_ _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4471_ as2650.r123\[1\]\[7\] as2650.r123\[0\]\[7\] as2650.r123_2\[1\]\[7\] as2650.r123_2\[0\]\[7\]
+ _4060_ _4064_ _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7700__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8963__CLK clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ net46 _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7190_ _2458_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _1493_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8256__A2 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _1290_ _1438_ _1441_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _4280_ _4285_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4509__I _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6724__I _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6974_ _2281_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8144__C _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8713_ _3884_ _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8644_ _1436_ _1782_ _1783_ _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_80_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _4279_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8192__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4807_ _4400_ _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8575_ _2410_ _3415_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8160__B _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5787_ as2650.holding_reg\[7\] _4397_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7526_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4738_ _4264_ as2650.cycle\[3\] _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7457_ _2712_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ net6 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6408_ _1691_ _1741_ _1742_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7388_ _2641_ _2644_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9127_ _0224_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6339_ _0883_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7290__I _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6258__A1 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9058_ _0155_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8798__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8009_ _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__A1 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__B2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5233__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6981__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7465__I _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__A1 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8986__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7289__A3 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8238__A2 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8229__C _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7997__A1 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7997__B2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8245__B _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6544__I _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8410__A2 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6421__A1 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6972__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ _0817_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4983__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6690_ _2004_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7921__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8360_ _3422_ _3582_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5572_ _0820_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7311_ _4339_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ as2650.r0\[4\] _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8291_ _2536_ _3515_ _3516_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6488__A1 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7242_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9141__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _4047_ _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A1 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8229__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _2445_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_1__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ as2650.stack\[1\]\[13\] _1369_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7978__C _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _0313_ _0294_ _0427_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6660__A1 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8401__A2 _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6957_ _1089_ _2100_ _2265_ _2266_ _1836_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5908_ _1267_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8165__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6888_ _4198_ _1814_ _2200_ _2102_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5839_ _0744_ _1241_ _0577_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8627_ _2279_ _3834_ _3836_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7912__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4702__I _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8558_ _1212_ _3772_ _2402_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7509_ _0406_ _2739_ _2743_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8489_ _1752_ _1695_ _3696_ _3706_ _4368_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__A1 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8640__A2 _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8065__B _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__A2 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9014__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6954__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4965__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8156__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4568__I1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8459__A2 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7923__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5142__A1 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6890__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7860_ _0423_ _4402_ _4256_ _2486_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8395__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7198__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6811_ _2084_ _2085_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7791_ as2650.pc\[11\] _1657_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6945__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7993__I1 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6742_ _0807_ _2040_ _2056_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ _1985_ _1988_ _1989_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__8698__A2 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4522__I _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8412_ _1406_ _2999_ _3563_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ _0880_ _0783_ _1027_ _1029_ _0664_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8343_ _2366_ _2720_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5555_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5381__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4506_ _4099_ _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8274_ _1320_ _2788_ _3423_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5486_ _4143_ _0867_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7122__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7225_ _1253_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5133__A1 _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6881__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7156_ as2650.r123_2\[0\]\[2\] _2405_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _1459_ _1461_ _4329_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_112_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8664__I _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7087_ _1672_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6633__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6038_ as2650.r123\[0\]\[3\] _1373_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4495__I0 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6184__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__A1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7989_ _1276_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9187__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4947__A1 _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8138__A1 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8689__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8310__A1 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7113__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5124__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8074__B1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8613__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7411__C _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__B _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A1 _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8523__B _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__A1 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5866__C _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8129__A1 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ as2650.holding_reg\[1\] _4376_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8301__A1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8301__B2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5115__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5271_ _0560_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7655__A3 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7010_ _2037_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7407__A3 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8604__A2 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7321__C _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8961_ _0072_ clknet_3_5__leaf_wb_clk_i as2650.r123_2\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7912_ _2380_ _2478_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8368__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8892_ _1654_ _1461_ _1470_ _4036_ _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_52_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4641__A3 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7843_ _2768_ _3070_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7040__A1 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7774_ _3015_ _3023_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4986_ _4414_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6725_ _1835_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6656_ _4108_ _1182_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7343__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8540__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _4124_ _0945_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5354__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _1901_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5538_ _4177_ _4178_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8326_ _1511_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8257_ _3175_ _3477_ _3483_ _3455_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5083__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8843__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7208_ _0812_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8188_ _4361_ _3405_ _2548_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _1852_ _2406_ _2413_ _2415_ _2416_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5811__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7231__C _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4880__A3 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__B _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7738__I _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5258__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8531__A1 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5345__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5896__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__B _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8598__A1 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A2 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5820__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6552__I _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4840_ as2650.cycle\[5\] _4433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7573__A2 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8770__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5584__A1 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _4364_ _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6510_ _1811_ _1814_ _1822_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_7490_ _2736_ _2679_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__A3 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8522__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _1770_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7876__A3 _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9160_ _0257_ clknet_leaf_71_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7316__C _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8111_ _3334_ _3338_ _3341_ _0424_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5323_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9091_ _0188_ clknet_leaf_9_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8042_ _1287_ _1275_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5639__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5254_ _0545_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6727__I _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ _0591_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8589__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8589__B2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7261__A1 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8944_ _0055_ clknet_leaf_51_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8875_ _3174_ _2377_ _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__I _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ _3070_ _3073_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6367__A3 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4969_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7757_ _2371_ _3005_ _3006_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _4138_ _1859_ _4091_ _4149_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7688_ _2936_ _2939_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7316__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7507__B _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7293__I _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6639_ _1862_ _1951_ _1955_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7867__A3 _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5878__A2 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8309_ _2879_ _3513_ _1380_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8277__B1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8816__A2 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4605__A3 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__A1 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7004__B2 as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6372__I _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8201__B1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8752__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7858__A3 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__I _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8807__A2 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7491__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8762__I _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7243__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7243__B2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6990_ _2291_ _2292_ _2294_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5941_ _1333_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5872_ as2650.pc\[0\] _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8660_ _1798_ _3849_ _3856_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8743__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7611_ _2601_ _1673_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4823_ _4410_ _4413_ _4416_ _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8591_ _1640_ _3803_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4754_ _4347_ _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7542_ _1020_ _1034_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7473_ _1298_ _2533_ _2727_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4685_ _4278_ _4240_ _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8002__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6424_ _0342_ _1677_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6355_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9143_ _0240_ clknet_leaf_37_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5306_ as2650.stack\[5\]\[8\] _0705_ _0711_ as2650.stack\[4\]\[8\] as2650.stack\[7\]\[8\]
+ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_9074_ _0171_ clknet_leaf_18_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6286_ _1622_ _1496_ _1520_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_88_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6457__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5237_ as2650.idx_ctrl\[0\] _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8025_ _3257_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5361__I _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7234__A1 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5099_ _0511_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8927_ _0038_ clknet_leaf_36_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8858_ _1491_ _3987_ _3995_ _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7537__A2 _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8734__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7809_ _3049_ _2542_ _3057_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5548__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8789_ _0383_ _0442_ _3370_ _0388_ _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8621__B _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_70_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8068__B _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7473__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__A3 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7473__B2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7776__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5787__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4615__I _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5539__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7926__I _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6830__I _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _4063_ _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7700__A2 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5711__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ as2650.stack\[0\]\[1\] _1439_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5181__I _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5022_ _4281_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A3 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8425__C _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9070__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8712_ as2650.r123\[1\]\[1\] _3890_ _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5924_ as2650.pc\[6\] _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8177__C1 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8643_ _2299_ _3840_ _3845_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5855_ _1245_ _1251_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8192__A2 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ _4388_ _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8574_ as2650.psu\[4\] _3772_ _1460_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5786_ _1187_ _0640_ _1188_ _4379_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_119_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7525_ _2528_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4753__A2 as2650.cycle\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ _4292_ _4312_ _4321_ _4330_ _4331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_108_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _0425_ _0357_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4668_ _4261_ _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _1619_ _0373_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7387_ _2641_ _2644_ _0641_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4599_ _4176_ _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9126_ _0223_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _0787_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6187__I _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9057_ _0154_ clknet_leaf_70_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6269_ as2650.psl\[1\] _1195_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5466__B1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8008_ _2454_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8616__B _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7947__S _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8707__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A2 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8183__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7930__A2 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4744__A2 _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5266__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7694__A1 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9093__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7430__B _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6421__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4983__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8174__A2 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8930__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6185__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _0721_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5571_ _0972_ _0974_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_129_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7310_ _2568_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4522_ _4115_ _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _2554_ _3293_ _3501_ _2595_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6488__A2 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7241_ _4237_ _1278_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4453_ _4046_ _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5904__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7172_ as2650.r123_2\[0\]\[5\] _2437_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5160__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7437__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _0812_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5999__A1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8436__B _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _0424_ _0425_ _0298_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8155__C _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _1213_ _2102_ _1817_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7566__I _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ _1022_ _2049_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6470__I _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8626_ as2650.stack\[7\]\[0\] _3835_ _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5838_ _1240_ _0818_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7912__A2 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8557_ _3700_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5769_ _1161_ _1162_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7508_ _2753_ _2763_ _4336_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8488_ _1695_ _1651_ _3705_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7676__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ net31 net30 net29 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5814__I _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5151__A2 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9109_ _0206_ clknet_leaf_27_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8953__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__A2 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8156__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__I _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4568__I2 as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7419__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8092__A1 _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6555__I _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__A1 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6810_ _2080_ _2083_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7790_ _2526_ _3037_ _3039_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6741_ _1850_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8147__A2 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4803__I _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__A1 _4439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6672_ as2650.r0\[2\] _1858_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8411_ _4425_ _3629_ _3631_ _3162_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5623_ _1028_ _0794_ _0548_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8342_ _0410_ _2984_ _3565_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5381__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5554_ _4207_ _0959_ _0943_ _0655_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _4098_ _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8273_ _3391_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5485_ _0892_ _0870_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7224_ _1635_ _2479_ _0339_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5133__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6330__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8607__B1 _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6881__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7155_ _2111_ _2419_ _2420_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8083__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6106_ _4047_ _0738_ _0485_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7086_ _2373_ _2360_ _2375_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7830__A1 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6633__A2 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8976__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _1392_ _1410_ _1411_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4495__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__A2 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7988_ _2781_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8613__C _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6939_ _2225_ _2248_ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4947__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8138__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5809__I _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__B2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7897__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8609_ _4188_ _0466_ _3812_ _3820_ _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7649__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5544__I _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8310__A2 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5124__A2 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8074__B2 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__I _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8804__B _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9131__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4938__A2 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__A1 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7888__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7934__I _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8301__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _4393_ _0678_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6312__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__A2 as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8065__A1 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7812__A1 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8960_ _0071_ clknet_leaf_75_wb_clk_i as2650.r123_2\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4626__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7911_ _1482_ _3153_ _3154_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_110_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8891_ _0494_ _0666_ _4398_ _4025_ _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7842_ net53 _2542_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7040__A2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7773_ _3017_ _3022_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4985_ _4350_ _0303_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5629__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8005__I _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6724_ _1833_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7879__A1 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6655_ _4061_ as2650.r123_2\[0\]\[7\] _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8540__A2 _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5606_ _4174_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5354__A2 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _0844_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8325_ _0395_ _3536_ _3549_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5537_ _0941_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8256_ _3260_ _3462_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6303__A1 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ _0844_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9004__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7207_ _0451_ _2340_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8675__I _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8187_ _4049_ _3395_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5399_ _0544_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7138_ _2404_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7803__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4708__I as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7069_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9154__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 as2650.cycle\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7955__S _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5593__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6790__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5345__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7885__A4 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8295__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8047__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8598__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8253__C _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7022__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4770_ _4311_ _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6128__A4 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5336__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__B1 _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6371_ net10 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8110_ _3339_ _3326_ _3340_ _0415_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5322_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9090_ _0187_ clknet_leaf_9_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8041_ _3263_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9177__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5184_ _0586_ _0592_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8943_ _0054_ clknet_leaf_50_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8874_ _3202_ _4022_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8163__C _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8210__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7825_ _3045_ _3003_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5024__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5024__B2 _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7756_ _2920_ _2921_ _3002_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4968_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ as2650.r0\[2\] _4090_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7574__I _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7687_ _2858_ _2937_ _2938_ _2882_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4899_ _0322_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _1952_ _1953_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6524__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A3 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _1881_ _1883_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8308_ _1379_ as2650.pc\[7\] _3513_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8277__A1 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8277__B2 as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8239_ _1092_ _4111_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8029__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7252__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8354__B _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5263__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A4 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8073__C _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7004__A2 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8752__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7484__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__A4 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7491__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7243__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8440__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _1267_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7610_ _2863_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4822_ _4415_ _4409_ _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8590_ _3800_ _3801_ _3802_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7541_ _1490_ _2760_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4753_ _4263_ as2650.cycle\[11\] _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5907__I _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7472_ _2728_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4684_ _4232_ _4250_ _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _1751_ _1753_ _1759_ _4372_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9142_ _0239_ clknet_leaf_37_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6354_ _4414_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5305_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9073_ _0170_ clknet_leaf_17_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6285_ _0487_ _1623_ _1462_ _4371_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8158__C _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8024_ _4301_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5236_ _0645_ _0597_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7997__C _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5167_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8431__A1 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ as2650.r123\[3\]\[5\] _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6473__I _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8926_ _0037_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6993__A1 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8857_ _3202_ _4007_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8902__B _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8734__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7808_ _2537_ _3056_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8788_ _4424_ _3515_ _3941_ _4436_ _4301_ _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5548__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7739_ _2553_ _2980_ _2988_ _2989_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8498__A1 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7170__A1 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7170__B2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5720__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7473__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8422__A1 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A2 _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5727__I _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7161__A1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7700__A3 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6558__I _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _1284_ _1438_ _1440_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8413__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A4 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4806__I _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6972_ _2280_ _0711_ _1270_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5778__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8711_ _3887_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5923_ _1121_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8177__B1 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8177__C2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8642_ as2650.stack\[7\]\[7\] _3841_ _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5854_ _4243_ _0462_ _1253_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_62_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _4388_ _4391_ _4392_ _4398_ _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_8573_ _0555_ _3738_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5785_ _0670_ _0640_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7524_ _2767_ _2534_ _2779_ _2729_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8013__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4736_ _4311_ _4262_ _4323_ _4329_ _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7455_ _0434_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4667_ _4260_ _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _1614_ _1737_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4697__B _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7386_ _2642_ _2643_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5702__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _4191_ _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9125_ _0222_ clknet_leaf_34_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6337_ _0676_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8652__A1 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9056_ _0153_ clknet_leaf_44_wb_clk_i as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6268_ _1596_ _1602_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8007_ _3235_ _3237_ _3239_ _1277_ _3033_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5219_ _0592_ _0593_ _0605_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6199_ _0880_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8404__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8909_ _0020_ clknet_leaf_75_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8707__A2 _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A3 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8351__C _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4451__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7694__A2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8891__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__I _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8643__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5457__A1 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__C _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6957__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8159__B1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__A3 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ as2650.stack\[6\]\[11\] _0719_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _4107_ _4112_ _4114_ _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7134__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7240_ _0471_ _1266_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8882__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ _4045_ _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6488__A3 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _2222_ _2406_ _2416_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5160__A3 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _0445_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A1 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7621__B _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ as2650.r123\[0\]\[5\] _1374_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5920__I _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5004_ _0365_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8008__I _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6955_ _1217_ _1840_ _2264_ _1810_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_74_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5906_ as2650.pc\[4\] _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_74_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6886_ _1009_ _2059_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8625_ _3833_ _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5837_ _1211_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7373__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5367__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8556_ as2650.psu\[3\] _3738_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5768_ _1004_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7507_ _2758_ _2761_ _2762_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _4261_ _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7125__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8487_ _0489_ _3256_ _3704_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5699_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7438_ _2684_ _2687_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8873__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7369_ _2592_ _2525_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9108_ _0205_ clknet_leaf_25_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5439__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9039_ _0007_ clknet_leaf_13_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6167__A2 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4568__I3 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8864__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9060__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8616__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8092__A2 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__S _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__A2 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A1 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _0802_ _2041_ _1834_ _2055_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ as2650.r0\[3\] _1860_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5187__I as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8410_ _2378_ _2722_ _3630_ _3139_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5622_ _4202_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__B1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8341_ _2965_ _0391_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ _0945_ _0799_ _0946_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5915__I _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ as2650.r0\[6\] _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8272_ _0335_ _3498_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8855__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5484_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5669__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ net24 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5133__A3 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6330__A2 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7154_ _2421_ _2422_ _2423_ _1545_ _2429_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8607__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8607__B2 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8447__B _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _0731_ _0501_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7085_ _2374_ _2367_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5650__I _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ as2650.r123_2\[0\]\[3\] _1391_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7830__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7987_ _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _2223_ _2235_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _4099_ _4091_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6149__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8608_ _1659_ _3754_ _3755_ _3819_ _0426_ _1090_ _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_109_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9083__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8539_ _1640_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__I _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7649__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8846__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8074__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4635__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6388__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6391__I _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__A3 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5060__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7888__A2 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5735__I _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8837__A1 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6312__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5115__A3 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5470__I _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6076__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7812__A2 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__A2 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A1 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7910_ _2504_ _2512_ _2513_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8890_ _4034_ _4035_ _3647_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7841_ _2537_ _3088_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7576__A1 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ _2953_ _2966_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7040__A3 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4984_ _0333_ _4417_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6723_ _1832_ _1852_ _2039_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ _1881_ _1969_ _1970_ _1953_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_108_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _4133_ _0942_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6585_ _1890_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5354__A3 _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8324_ _3537_ _3532_ _3548_ _3188_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8021__I _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8828__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _4205_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8255_ _3282_ _3462_ _3481_ _3232_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8943__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7206_ _1526_ _2343_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8186_ _3411_ _3412_ _3413_ _3414_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4865__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8056__A2 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7137_ _1854_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ as2650.addr_buff\[0\] _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A2 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6019_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A1 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5042__A2 _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7319__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7319__B2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5555__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8819__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8295__A2 _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8047__A2 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5290__I _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7558__A1 _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8755__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__I as2650.alu_op\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7010__I _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8966__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__B2 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _0675_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5321_ _4380_ _0474_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6297__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8040_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5252_ _0601_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5183_ _0584_ _4395_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__A3 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8942_ _0053_ clknet_leaf_58_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8873_ as2650.overflow _4017_ _4021_ _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4544__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7824_ _3070_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8210__A2 _4448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5024__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7755_ _2971_ _2975_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4967_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6772__A2 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6706_ _1969_ _2020_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7686_ as2650.pc\[7\] _1141_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4898_ _0324_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _4105_ _1895_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5375__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _1879_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8307_ _3531_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5519_ _0771_ _0767_ _0848_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__8686__I _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8277__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6499_ _4393_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6288__A1 _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8619__C _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8238_ _1092_ _4111_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__I _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8169_ _3362_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4454__I _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8201__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8989__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7960__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7712__A1 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5723__B1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6279__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7779__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8440__A2 _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8728__B1 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5870_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5006__A2 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4821_ _4414_ _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7951__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7540_ _0314_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4752_ _4345_ _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ _2532_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _4268_ _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6506__A2 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _1758_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9144__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9141_ _0238_ clknet_leaf_37_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5190__A1 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _4402_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5923__I _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9072_ _0169_ clknet_leaf_17_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6284_ _4329_ _1459_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8023_ _0973_ _3249_ _3253_ _3255_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5235_ _0596_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5166_ _4259_ _0571_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_84_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8455__B _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5097_ _0510_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8925_ _0036_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8856_ _0610_ _3996_ _4000_ _4006_ _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8195__A1 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7807_ _3040_ _3055_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8787_ _0460_ _2336_ _0389_ _0360_ _0490_ _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_5999_ as2650.r123_2\[0\]\[0\] _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4756__A1 _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7518__C _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ _2330_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ _2263_ _1233_ _0640_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4508__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5236__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__B2 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9017__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6984__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4912__I _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8489__A2 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A1 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__A1 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__A2 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5020_ _0357_ _4442_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6672__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8413__A2 _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _1366_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6975__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8710_ _0696_ _3883_ _3889_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _1302_ _1317_ _1318_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8177__A1 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8177__B2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7619__B _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5853_ _0614_ _0359_ _1245_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_62_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8641_ _2297_ _3840_ _3844_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7924__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4804_ _4393_ _4397_ _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_72_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5784_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8572_ _3691_ _1009_ _3784_ _3785_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _2772_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _4328_ _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7454_ net55 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ net6 as2650.cycle\[13\] _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _1474_ _0371_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5163__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ _0883_ _0896_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4597_ _4190_ _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9124_ _0221_ clknet_leaf_81_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6336_ _1672_ _1095_ _1674_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8101__A1 _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9055_ _0152_ clknet_leaf_45_wb_clk_i as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6267_ _1191_ _1185_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8652__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8006_ _3238_ _2331_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5218_ _0581_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _1530_ _1547_ _1548_ _1549_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8404__A2 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _4310_ _0556_ _0557_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_84_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6966__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__A1 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8908_ _0019_ clknet_leaf_66_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8168__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7529__B _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8839_ _1625_ _1641_ _1634_ _3989_ _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7915__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6718__A2 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A4 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8340__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5154__A1 _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5563__I _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8891__A2 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8079__C _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6654__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4907__I _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8159__A1 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6343__B _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7382__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4520_ _4068_ _4113_ _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8331__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4451_ as2650.cycle\[6\] _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5473__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6893__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5696__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7170_ _2037_ _2414_ _2411_ _1312_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5160__A4 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _1131_ _1469_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5448__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _1392_ _1423_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _4324_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8398__A1 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6954_ _2263_ _1840_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5905_ _1018_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6885_ _2195_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8024__I _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8624_ _3833_ _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5836_ _1133_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_50_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8570__A1 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5767_ _1165_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8555_ _1701_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7506_ _0326_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4718_ _4301_ _4308_ _4311_ _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8322__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7125__A2 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8486_ _3699_ _3702_ _3703_ _1700_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5698_ _1055_ _0959_ _1081_ _1032_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_120_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8322__B2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A1 _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7437_ _2373_ _2564_ _2692_ _2693_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4649_ as2650.halted _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8873__A2 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _2582_ _2583_ _2626_ _0458_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9107_ _0204_ clknet_leaf_24_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6319_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7299_ _2547_ _2558_ _4242_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6636__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5439__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9038_ _0006_ clknet_leaf_14_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7103__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8313__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7116__A2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8818__B _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8616__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8537__C _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _1984_ _1985_ _1986_ _1949_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1023_ _0788_ _1025_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5366__B2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8340_ _1390_ _3533_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5552_ _0658_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8304__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4503_ _4072_ _4096_ _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8271_ _1322_ _3269_ _3497_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5483_ _0645_ _0597_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8855__A2 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6866__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5669__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7222_ _4392_ _2481_ _2483_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7153_ _0908_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8607__A2 _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _0562_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7084_ as2650.addr_buff\[3\] _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _1409_ _1382_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8019__I _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7986_ _3216_ _3218_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8791__A1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _2223_ _2235_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__I _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _2161_ _2163_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_74_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7346__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8607_ _1028_ _3777_ _3695_ _1619_ _3818_ _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5819_ _1211_ _0878_ _0661_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _2063_ _2093_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8538_ _0454_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__A2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8846__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8469_ _3686_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6609__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4457__I _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7034__A1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8782__A1 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5596__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5288__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7888__A3 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__A3 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8837__A2 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5115__A4 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7273__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5823__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7840_ _3084_ _3087_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8773__A1 as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7771_ _0418_ _3020_ _2943_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _0318_ _0406_ _0330_ _0328_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ as2650.r123_2\[2\]\[0\] _1856_ _2036_ _2038_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8525__A1 _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6653_ _4128_ _1874_ _1872_ _1968_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5926__I _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6531__B _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__I _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _0804_ _0891_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_118_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _1876_ _1897_ _1899_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8323_ _4429_ _3542_ _3547_ _3139_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_121_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5535_ _4136_ _4141_ _4147_ _4153_ _0798_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_106_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8828__A2 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8254_ _3473_ _3474_ _3480_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5466_ _0655_ _0868_ _0870_ _0871_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__6303__A3 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8458__B _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7205_ _2460_ _1434_ _2468_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8185_ as2650.stack\[5\]\[4\] _2455_ _3379_ as2650.stack\[4\]\[4\] _0905_ _3414_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_82_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5397_ _4208_ _0798_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7136_ _2402_ _1815_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8056__A3 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7067_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ as2650.r123\[0\]\[1\] _1373_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8764__A1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A1 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9050__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7969_ as2650.psu\[7\] _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7319__A2 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__A1 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8819__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8368__B _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_33_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5502__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__A1 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7007__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__B _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7558__A2 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__A1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7730__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ _0716_ _0724_ _0729_ _0723_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _0537_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6297__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5182_ _4164_ _0587_ _0590_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_68_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A1 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8941_ _0052_ clknet_leaf_58_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9073__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__I _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8872_ _0387_ _4018_ _4017_ _4020_ _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4480__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8746__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7823_ _3045_ _3006_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__A2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7754_ _2371_ _3001_ _3003_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4966_ net3 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6705_ _1954_ _2021_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7685_ _2853_ _2881_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_71_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4897_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4560__I _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6636_ as2650.r0\[6\] _1868_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5732__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__A2 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _1880_ _1881_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_106_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8306_ _1379_ _3530_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7804__C _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5518_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8188__B _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6498_ _4356_ _1807_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7485__A1 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6288__A2 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6487__I _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8237_ _1657_ _4096_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5449_ _0624_ _0848_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5496__B1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8168_ _1305_ _3396_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _1796_ _2393_ _2399_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8099_ _2713_ _3326_ _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7960__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5971__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5566__I _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4470__I _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7476__A1 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6279__A2 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9096__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7228__A1 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7779__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8545__C _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6451__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4645__I _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8728__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4462__A1 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8728__B2 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6203__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7400__A1 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8933__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ net3 _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7951__A2 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4751_ _4344_ _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7470_ _2719_ _2726_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4682_ _4254_ _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8900__A1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6421_ _1754_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7691__I _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9140_ _0237_ clknet_leaf_37_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6352_ as2650.psl\[7\] _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7467__A1 _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9071_ _0168_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6283_ _0552_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8022_ as2650.stack\[4\]\[0\] _3254_ _0906_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7219__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7640__B _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _0547_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ as2650.r123\[3\]\[4\] _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8431__A3 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8027__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6442__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8924_ _0035_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8855_ _2961_ _0914_ _4005_ _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8195__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7806_ _3015_ _3023_ _3041_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8786_ _1479_ _2639_ _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7737_ _2978_ _4431_ _2721_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4756__A2 _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5953__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _0369_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ _1215_ _1233_ _2899_ _2900_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _1893_ _1908_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7599_ as2650.pc\[6\] _1656_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A1 _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8365__C _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__I _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6433__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8956__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5944__A1 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8400__I _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5172__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__A2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__A1 _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6970_ _1283_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ as2650.stack\[3\]\[5\] _1310_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8177__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8640_ as2650.stack\[7\]\[6\] _3841_ _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5852_ _0460_ _1249_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9111__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7924__A2 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _4396_ _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4738__A2 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5935__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8571_ _3765_ _1015_ _3686_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5783_ _4076_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7522_ _2740_ _0393_ _2714_ _2777_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4734_ _4325_ _4327_ _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7688__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7453_ as2650.pc\[3\] _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ net5 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6404_ _1590_ _1208_ _1610_ _4050_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7354__C _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7384_ _0893_ _0895_ _1717_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5163__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _4136_ _4141_ _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9123_ _0220_ clknet_leaf_82_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6335_ _1673_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8101__A2 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9054_ _0151_ clknet_leaf_46_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6112__A1 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6266_ _1201_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8466__B _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _3128_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7860__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8979__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _0605_ _0592_ _0593_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6197_ _0469_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8185__C _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _4057_ _0492_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7612__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5079_ _0485_ _0487_ _0489_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_44_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8907_ _0018_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4977__A2 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8838_ _0454_ _0364_ _1515_ _3988_ _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_44_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7915__A2 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8769_ as2650.stack\[4\]\[3\] _3926_ _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__I as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5154__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7851__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6406__A2 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8159__A2 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4923__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7906__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6590__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8331__A2 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6342__A1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8619__B1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__A1 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6120_ _0739_ _1472_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5448__A3 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7842__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ as2650.r123_2\[0\]\[5\] _1376_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5853__B1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5002_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _1214_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A1 _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5929__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ _1271_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6884_ _2173_ _2196_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8623_ _1346_ _1349_ _1351_ _1347_ _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5835_ _0748_ _1209_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8570__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8554_ _1589_ _3768_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5766_ _1069_ _1067_ _1070_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7365__B _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7505_ _2376_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4717_ _4310_ _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8485_ _1923_ _1472_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5697_ _1082_ _1083_ _0871_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__8322__A2 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8040__I _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _2345_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4648_ _4241_ _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7367_ _1288_ _0380_ _2605_ _2606_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_2_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4579_ _4172_ _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9106_ _0203_ clknet_leaf_25_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8086__A1 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6318_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7812__C _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7298_ _2541_ _4437_ _2549_ _2557_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7833__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9037_ _0005_ clknet_leaf_13_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6636__A2 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6249_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9157__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8546__C1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8010__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8313__A2 _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A1 _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__A1 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7722__C _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7824__A1 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A2 _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A1 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8001__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8552__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5620_ _0521_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6563__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _0949_ _0878_ _0661_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _4063_ _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5118__A2 _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8270_ _3273_ _3462_ _3486_ _3496_ _3313_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5417__C _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _0652_ _0875_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7221_ net23 _2481_ _2482_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6866__A2 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4877__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8068__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6330__A4 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7152_ _2408_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7815__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ as2650.psu\[5\] _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4828__I _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7815__B2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _1710_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8463__C _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7985_ _2519_ _3217_ _3101_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5054__A1 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__I as2650.alu_op\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8791__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _1177_ _2246_ _2096_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6867_ _1087_ _2156_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8606_ _3813_ _3817_ _0448_ _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ _1089_ _0669_ _1220_ _0689_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5357__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6798_ _2065_ _2092_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8537_ _0355_ _1591_ _3751_ _3752_ _3693_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_109_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5749_ _4181_ _1010_ _1134_ _0941_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_108_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A2 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6306__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _4282_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4580__A3 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7419_ _1689_ _2674_ _2676_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_135_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6857__A2 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8399_ _3316_ _3604_ _3617_ _3620_ _3220_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8059__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6953__I _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__A1 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7034__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6174__B _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8782__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7888__A4 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8298__A1 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8829__B _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__A1 _4448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__B _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__I _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8222__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5036__A1 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7770_ _3015_ _3019_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4982_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6721_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _1968_ _1875_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6536__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4547__B1 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6583_ _0588_ _1882_ _1896_ _4139_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8322_ _2531_ _3531_ _3544_ _0358_ _3546_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8289__A1 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__I as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _0804_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8253_ _2531_ _3461_ _3478_ _3479_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _4143_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7204_ as2650.stack\[2\]\[14\] _2458_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8184_ as2650.stack\[7\]\[4\] _2388_ _3347_ as2650.stack\[6\]\[4\] _3413_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _4176_ _0804_ _0648_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7135_ _0730_ _2409_ _2412_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8461__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7066_ _2358_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _1390_ _1391_ _1392_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__C _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__I _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A2 _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7968_ _0336_ _3201_ _3202_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7818__B _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6919_ _1120_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7899_ net52 _0299_ _0380_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8516__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__B1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8819__A3 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_73_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8452__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7007__A2 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8204__B2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8755__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8507__A2 _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_3_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8278__C _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5250_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5181_ _4375_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7246__A2 _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8443__A1 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5257__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8940_ _0051_ clknet_leaf_58_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6526__C _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8871_ _1691_ _3182_ _4019_ _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5009__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8746__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4480__A2 _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7822_ as2650.addr_buff\[4\] _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5002__I _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7753_ _2907_ _2924_ _2926_ _3002_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4965_ _0388_ _4314_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6704_ _4075_ _1882_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ as2650.pc\[8\] _1140_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4896_ _4412_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5158__B _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6635_ _4127_ _1874_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _4150_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8305_ _1327_ _3500_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5517_ _0922_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6497_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8236_ _2355_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _4251_ _0631_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6288__A3 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8167_ _1297_ _3359_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5379_ _0682_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7118_ as2650.stack\[4\]\[12\] _2395_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8434__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8098_ _2369_ _3292_ _3327_ _2596_ _3328_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ _4256_ _4287_ _0552_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6996__A1 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6008__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4751__I _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5723__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5582__I _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8673__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__C _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__A1 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__B1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__B1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8842__B _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4462__A2 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8728__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7400__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4750_ net6 as2650.cycle\[13\] _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4681_ _4270_ _4272_ _4274_ _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7164__A1 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ _0339_ _4246_ _4256_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__8900__A2 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7905__C _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A2 _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6588__I _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ _1686_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ as2650.psu\[0\] as2650.psu\[1\] _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7467__A2 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9070_ _0167_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6282_ _0373_ _1618_ _1620_ _1225_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5478__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9040__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8021_ _3244_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5233_ _0318_ _0526_ _0528_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_97_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A2 _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8416__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _0509_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9190__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8923_ _0034_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8854_ _0931_ _4003_ _4004_ _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7805_ _0418_ _3043_ _3053_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8785_ _3378_ _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5997_ _0549_ _1280_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8043__I _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__I _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7736_ _2550_ _2970_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4948_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__A3 _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7667_ _2787_ _2918_ _2919_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7155__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4879_ _4433_ _4283_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7882__I _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _1921_ _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7598_ _0405_ _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6902__A1 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ _4160_ _1864_ _1865_ _0752_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8219_ _1019_ _4120_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8407__A1 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A2 _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__A1 _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5492__I1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7993__S _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4481__I as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5944__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8894__A1 _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9063__CLK clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8128__I _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _0341_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_94_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7385__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ _4395_ _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8570_ _2762_ _1035_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5782_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _1693_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4733_ _4306_ _4326_ _4327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7137__A1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7452_ _2699_ _2708_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8885__A1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ _4051_ _4222_ _4237_ _4257_ _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_6403_ _1694_ _1695_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7383_ _2569_ _2615_ _2640_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4595_ _4126_ _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9122_ _0219_ clknet_leaf_81_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6334_ _1143_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8637__A1 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9053_ _0150_ clknet_leaf_53_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6265_ _1164_ _1603_ _1595_ _1073_ _1202_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5950__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6112__A2 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8004_ _1676_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5216_ _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6196_ net44 _1538_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7860__A2 _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4566__I _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _4046_ _4438_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7612__A2 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5078_ _0305_ _0490_ _0491_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_85_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5623__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6781__I _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8906_ _0017_ clknet_leaf_60_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8837_ _4251_ _2343_ _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8768_ _2287_ _3925_ _3929_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7719_ as2650.addr_buff\[1\] _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8699_ as2650.stack\[5\]\[13\] _3872_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8876__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8628__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7300__A1 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8923__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7064__B1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7603__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8800__A1 _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8392__B _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6905__B _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7367__B2 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7119__A1 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6590__A2 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8867__A1 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8619__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8619__B2 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__B _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8095__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1422_ _1382_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7842__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input7_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5853__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A2 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _4367_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _1831_ _2247_ _2262_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A2 _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _1272_ _1300_ _1301_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6883_ _2114_ _2140_ _2172_ _2175_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _0580_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8622_ _3825_ _3831_ _3832_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__A1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5765_ _1165_ _1167_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8553_ _3691_ _0940_ _3767_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7504_ _2759_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4592__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ _4309_ _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8484_ _0610_ _3701_ _0574_ _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8858__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5696_ _1088_ _0779_ _1098_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7435_ _2564_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4647_ _4240_ _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8946__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _2607_ _2621_ _2623_ _2624_ _2574_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4578_ _4107_ _4112_ _4114_ _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_89_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9105_ _0202_ clknet_leaf_25_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6317_ net2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8086__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7297_ _2540_ _2551_ _2553_ _2556_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9036_ _0000_ clknet_leaf_18_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6248_ _1513_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _1532_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7597__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_3_0_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8794__B1 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8546__B1 _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8546__C2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_27_wb_clk_i clknet_3_6__leaf_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4583__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8849__A1 _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6324__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__A3 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7521__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6686__I _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8077__A2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__I _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__I _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5063__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4810__A2 _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8001__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8969__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7760__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _0950_ _0879_ _0956_ _0689_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4574__A1 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _4083_ _4087_ _4092_ _4094_ _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _0877_ _0878_ _0661_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5118__A3 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _1686_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8297__B _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4877__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7151_ _2427_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8068__A2 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1457_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7815__A2 _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7082_ _2369_ _2360_ _2372_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A2 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5826__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6033_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7579__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4844__I _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8240__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7220__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7984_ _2768_ _4241_ _2863_ _4286_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5054__A2 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _1154_ _2040_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _2168_ _2170_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8605_ _4092_ _1472_ _2402_ _3816_ _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5817_ _1026_ _1213_ _1219_ _0879_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6797_ _1855_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8536_ _3688_ _0896_ _0354_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5748_ _0648_ _1135_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__A1 _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6306__A2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ _1082_ _1083_ _0892_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8467_ _3684_ _3685_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7418_ _2630_ _2675_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_136_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8398_ _3606_ _3618_ _3619_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8059__A2 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _0785_ _0801_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8000__B _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9019_ _0130_ clknet_leaf_31_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6490__A1 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8231__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5596__A3 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7990__A1 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A2 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8298__A2 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4859__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4929__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8222__A2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4981_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8580__B _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7981__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6720_ _1853_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ as2650.r0\[5\] _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6536__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ _0636_ _0986_ _1001_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4547__A1 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _4128_ _1898_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9147__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8321_ _0411_ _2955_ _3545_ _3475_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5533_ _0914_ _0916_ _0929_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8289__A2 _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8252_ _1143_ _0463_ _3370_ _2382_ _4360_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5464_ _0654_ _0657_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7203_ _2460_ _1427_ _2467_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4839__I _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8183_ as2650.stack\[1\]\[4\] _3252_ _3379_ as2650.stack\[0\]\[4\] _1046_ _3412_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5395_ as2650.idx_ctrl\[1\] _0647_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7134_ _0663_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7065_ _2333_ _2339_ _2351_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6016_ as2650.r123_2\[0\]\[1\] _1376_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6472__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8046__I _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5027__A2 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8490__B _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7967_ _0469_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7972__A1 _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4786__A1 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6918_ _2156_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7898_ _2385_ _0415_ _3143_ _0438_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7724__A1 _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6849_ _2129_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6527__A2 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8519_ _0355_ _0775_ _3733_ _3735_ _3693_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8384__C _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7795__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A1 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6204__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7191__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8691__A2 _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7035__I _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6__f_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _0589_ _0539_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A3 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8443__A2 _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__A2 _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8870_ _1732_ _3180_ _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5009__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7821_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7752_ as2650.addr_buff\[0\] as2650.addr_buff\[1\] as2650.addr_buff\[2\] _3002_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4964_ _0359_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _4075_ _1895_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7683_ _2795_ _2930_ _2934_ _2700_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4895_ _0323_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6634_ _1948_ _1949_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5193__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _1875_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8304_ _1328_ _3499_ _3528_ _3529_ _0334_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5516_ _0916_ _0921_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6496_ _0553_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8131__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8235_ _3461_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5447_ _4389_ _4299_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8682__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8166_ _3394_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5378_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7117_ _1794_ _2392_ _2398_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8097_ as2650.addr_buff\[2\] _3140_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8434__A2 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5248__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7048_ _1518_ _2340_ _0434_ _1514_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4551__S0 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8999_ _0110_ clknet_leaf_52_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7945__A1 _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__B1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8370__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6381__B1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8379__C _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6684__A1 _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6908__B _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7228__A3 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8425__A2 _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5239__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__B2 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5531__C _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4998__B2 _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4942__I _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4680_ _4273_ as2650.cycle\[5\] _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8361__A1 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6911__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6350_ _1685_ _1688_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6281_ _1619_ _0373_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5232_ _0314_ _0639_ _0641_ _0531_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__6675__A1 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8020_ as2650.stack\[7\]\[0\] _3250_ _3251_ as2650.stack\[6\]\[0\] _3252_ as2650.stack\[5\]\[0\]
+ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_88_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7219__A3 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5163_ _0488_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A1 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6427__B2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ as2650.r123\[3\]\[3\] _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6978__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8922_ _0033_ clknet_leaf_54_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5013__I _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8853_ _1192_ _1196_ _1200_ _1004_ _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__I _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ _2678_ _3048_ _3052_ _2620_ _0417_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8784_ _0321_ _1761_ _3938_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _1372_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5402__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7735_ _2978_ _2542_ _2985_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _4342_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ net54 _2829_ _2830_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4878_ _4271_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7384__B _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6617_ _1932_ _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5166__A1 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__I _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _2620_ _2850_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _1861_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8104__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8655__A2 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6479_ _1426_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6666__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8218_ _1019_ _4120_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7831__C _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6130__A3 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8407__A2 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8149_ _3243_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6418__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A3 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6969__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6019__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7918__A1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4762__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8343__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8894__A2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__A1 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7606__B1 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7082__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5632__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7909__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _4046_ _1246_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7385__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8582__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4801_ _4394_ _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A1 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _0671_ _1057_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _2773_ _2775_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4732_ _4269_ _4239_ _4157_ _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8334__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__A1 _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7451_ _2700_ _2706_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4663_ _4247_ _4256_ _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8885__A2 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6402_ _1699_ _1739_ _1639_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7382_ _0785_ _0806_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4594_ _4185_ _4187_ _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__8098__B1 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9121_ _0218_ clknet_leaf_81_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6333_ _1023_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5008__I _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6264_ _1062_ _1059_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9052_ _0149_ clknet_leaf_56_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8003_ _4161_ _2891_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5215_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__I _4439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5320__B2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _1545_ _1533_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7860__A3 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _0550_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8270__B1 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _0493_ _0496_ _4230_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5084__B1 _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6820__A1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8905_ _0016_ clknet_leaf_60_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4582__I _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8836_ _1614_ _3777_ _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8573__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8767_ as2650.stack\[4\]\[2\] _3926_ _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5979_ _1353_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7893__I _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7718_ _2966_ _2968_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8325__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8698_ _1796_ _3874_ _3880_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _1216_ _1234_ _2901_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8876__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6887__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7300__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7064__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8261__B1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4492__I _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7367__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8564__A1 _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8316__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7119__A2 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__I _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6212__I _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9180__CLK clknet_3_2__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6342__A3 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5550__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8619__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__I _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _4351_ _0421_ _0422_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5853__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7055__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8252__B1 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ as2650.r123_2\[2\]\[6\] _2112_ _2261_ _2142_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__I _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__A3 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5902_ as2650.stack\[3\]\[3\] _1285_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6882_ _2179_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8621_ _1240_ _3727_ _0351_ _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5833_ _1230_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8602__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8552_ _3765_ _0948_ _3766_ _3686_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5764_ _1165_ _1167_ _0930_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7503_ _4411_ _1531_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4715_ as2650.halted net5 _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8483_ _3700_ _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8858__A2 _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4592__A2 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5695_ _1099_ _0783_ _0779_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6869__A1 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7434_ _1679_ _0962_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4646_ _4238_ _4239_ _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7662__B _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ _2622_ _2589_ _0405_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4577_ _4169_ _4170_ _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_9104_ _0201_ clknet_leaf_27_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _0813_ _1468_ _0496_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7296_ _2555_ _2328_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9035_ _0146_ clknet_leaf_13_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6247_ _1578_ _1434_ _1586_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _0385_ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_97_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5129_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_73_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7597__A2 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8794__A1 _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8794__B2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8546__A1 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8546__B2 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8819_ _1463_ _2365_ _1496_ _3970_ _3971_ _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_3_5__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8512__I _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__A2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7128__I _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6032__I _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5532__A1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5871__I _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7588__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5599__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A3 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8537__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7760__A2 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7038__I _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ _4093_ _4085_ _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_118_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5480_ _0878_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ as2650.r123_2\[0\]\[1\] _2405_ _2426_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6101_ as2650.r123_2\[3\]\[7\] _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6079__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7081_ _2371_ _2367_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6032_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7579__A2 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8776__A1 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7983_ _3155_ _3213_ _3214_ _3215_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6117__I _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__A2 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _2238_ _2041_ _2097_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5021__I _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8528__A1 _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6865_ _1832_ _2153_ _2178_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8913__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8604_ _3814_ _3701_ _3815_ _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5816_ _1216_ _1024_ _1218_ _0685_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _0866_ _2096_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8535_ _3734_ _0874_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5747_ _0781_ _1138_ _1150_ _0899_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8466_ _1429_ _3622_ _3354_ _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5678_ _0951_ _4177_ _4178_ _4173_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7503__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8700__A1 _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7417_ _2523_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5514__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6787__I _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ as2650.psl\[7\] _4085_ _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8397_ _3487_ _0978_ _3551_ _3604_ _3495_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_85_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7348_ _0404_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5624__C _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8000__C _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _1276_ _2328_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5817__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9018_ _0129_ clknet_leaf_31_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6736__B _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8767__A1 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8519__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7990__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4770__I _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5753__A1 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9099__CLK clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4945__I _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6481__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6233__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8580__C _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6650_ _4105_ _1889_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ _0770_ _0996_ _1003_ _1004_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5744__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _1869_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8320_ _1380_ _2586_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5532_ _0931_ _0935_ _0936_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__8143__C1 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8251_ _3475_ _3477_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ _0657_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7202_ as2650.stack\[2\]\[13\] _2458_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8182_ as2650.stack\[3\]\[4\] _2388_ _3347_ as2650.stack\[2\]\[4\] _3411_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5394_ _0652_ _0802_ _0692_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7249__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7133_ _2410_ _1815_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8446__B1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5016__I _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _1488_ _0361_ _2354_ _2356_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4855__I _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _1371_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6472__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8749__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4483__A1 _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7966_ _4450_ _4399_ _1279_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7387__B _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _2227_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_78_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4786__A2 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5983__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__B _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7897_ net52 _3142_ _0414_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _2131_ _2132_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4538__A2 _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ as2650.r123_2\[2\]\[1\] _1856_ _2094_ _2038_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8518_ _3734_ _0802_ _0354_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8449_ _3648_ _3649_ _3668_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7406__I _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5499__B1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__A1 _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4765__I _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7412__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6980__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7963__A2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7297__B _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_82_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_82_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A4 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__A2 _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4529__A2 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7479__A1 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__I _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4675__I _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7651__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5257__A3 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7403__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7820_ as2650.pc\[12\] _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9114__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__B1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7751_ _2971_ _2973_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6702_ _1983_ _1991_ _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7682_ _2698_ _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4894_ _4273_ as2650.cycle\[3\] _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ as2650.r0\[0\] _4090_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6564_ _4127_ _1872_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6390__A1 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8303_ _3221_ _3502_ _3271_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5455__B _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5515_ _0916_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _0524_ _4310_ _0515_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8131__A2 _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8234_ _1321_ _3460_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5446_ _0850_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7890__A1 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ _2767_ _3393_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5377_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ as2650.stack\[4\]\[11\] _2395_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8096_ _2663_ _3317_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6286__B _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7642__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _1587_ _1519_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4551__S1 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8998_ _0109_ clknet_leaf_52_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5956__A1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7949_ _3170_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6381__B2 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__C _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7881__A1 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7228__A4 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6436__A2 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8189__A2 _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7739__C _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7936__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5947__A1 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8361__A2 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5300_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6280_ _4081_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5231_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4686__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _0477_ _0491_ _0482_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_68_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7624__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6427__A2 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5093_ _0508_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8921_ _0032_ clknet_leaf_35_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6834__B _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8852_ _4002_ _1596_ _1606_ _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7803_ _3049_ _3051_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_92_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8783_ _2377_ _1754_ _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7734_ _2903_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4946_ _4302_ _4055_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_71_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ _2879_ _2880_ _2917_ _0340_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4877_ _0298_ _0300_ _0304_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5964__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6616_ _1913_ _1917_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5166__A2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _2832_ _2849_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6547_ _1859_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8104__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6115__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _1796_ _1787_ _1797_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8496__B _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8217_ _3440_ _3444_ _3132_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5429_ as2650.holding_reg\[2\] _0602_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8148_ _3343_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A2 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4692__A4 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8079_ _1510_ _3275_ _3309_ _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__A2 _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5874__I _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6106__A1 _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7854__A1 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6657__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7606__A1 _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7606__B2 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8803__B1 _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5114__I _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8853__C _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7082__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7469__C _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8031__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ as2650.ins_reg\[3\] as2650.ins_reg\[2\] _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5780_ as2650.holding_reg\[7\] _1057_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _4324_ _4234_ _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5784__I _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8334__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7450_ _0338_ _2574_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4662_ _4255_ _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6345__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _1701_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6896__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7381_ _0883_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4593_ _4186_ _4168_ _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9120_ _0217_ clknet_leaf_80_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8098__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6332_ _0793_ _1213_ _1669_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7845__A1 _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6648__A2 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9051_ _0148_ clknet_leaf_54_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6263_ _0998_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7504__I _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8002_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5214_ _4390_ _0495_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6194_ _0950_ _1535_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7860__A4 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5145_ _0524_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__B1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__C2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8270__A1 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__A1 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__B2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__I _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8904_ _0015_ clknet_leaf_76_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8022__A1 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8835_ _3981_ _3985_ _3986_ _0349_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_4__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__A1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5387__A2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8766_ _2285_ _3925_ _3928_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5978_ _1353_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7781__B1 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7717_ _2967_ _2940_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8697_ as2650.stack\[5\]\[12\] _3876_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5694__I _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8070__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7648_ _2899_ _2900_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6336__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7579_ _1657_ _1137_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4898__A1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7836__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7064__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8261__A1 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8261__B2 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__I _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A1 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8564__A2 _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8316__A2 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6327__A1 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6342__A4 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7827__A1 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7827__B2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7324__I _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6368__C _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A2 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7055__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8252__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8252__B2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__A1 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4683__I _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6950_ _2250_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6802__A2 _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__A1 _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5901_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8004__A1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__A4 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6881_ _2190_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8620_ _1217_ _2606_ _3755_ _3829_ _3830_ _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _0899_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6566__A1 _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8551_ _2929_ _0962_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5763_ _1066_ _1074_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7502_ _2562_ _2757_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4714_ _4307_ _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8482_ _0480_ _0491_ _0478_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5694_ _4189_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7433_ _2650_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6869__A2 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4645_ _4052_ _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7364_ _2622_ _2589_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4576_ as2650.alu_op\[0\] as2650.alu_op\[1\] as2650.alu_op\[2\] _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9103_ _0200_ clknet_3_6__leaf_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7818__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _1465_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _2554_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9034_ _0145_ clknet_leaf_9_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6246_ as2650.stack\[3\]\[14\] _1576_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8491__A1 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__B1 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _0534_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8243__A1 _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7046__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5128_ _0529_ _0323_ _0525_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_85_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5057__A1 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8794__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8992__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _0477_ _4379_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_85_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9101__D _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8818_ _2410_ _3968_ _4361_ _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8749_ _0967_ _3906_ _3917_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5780__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__A3 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6324__A4 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7809__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4768__I _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__I _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8482__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_wb_clk_i clknet_3_7__leaf_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6983__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8234__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5599__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8537__A2 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8859__B _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6100_ _1456_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7080_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7989__I _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ as2650.pc\[11\] _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8225__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7028__A2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5039__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7982_ _3122_ _3125_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6251__A3 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6933_ _1121_ _2042_ _2043_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8528__A2 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ as2650.r123_2\[2\]\[3\] _2112_ _2177_ _2142_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7200__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8603_ _1660_ _3701_ _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5815_ _1217_ _0682_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6795_ _2057_ _2108_ _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__I _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8534_ _3730_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _1148_ _1149_ _0781_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8465_ _3316_ _3670_ _3680_ _3683_ _3271_ _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5677_ _4115_ _4125_ _0869_ _4199_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8700__A2 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7416_ _1292_ _2583_ _2672_ _2673_ _2525_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4628_ _4221_ _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8396_ _3176_ _3604_ _0436_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7347_ _4276_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _4152_ _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8464__A1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ _2537_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5278__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9017_ _0128_ clknet_leaf_30_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6229_ _1351_ _1574_ _1367_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8216__A1 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9170__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8519__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__B2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__I _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6702__A1 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4498__I _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__A1 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5269__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8207__A1 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8758__A2 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__I _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8391__B1 _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5600_ _0625_ _0992_ _0994_ _1005_ _0856_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6580_ _0588_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5531_ _0626_ _0922_ _0937_ _0632_ _0582_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_118_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8143__B1 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8143__C2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8250_ _1692_ _2869_ _3476_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8694__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _4190_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7201_ _2460_ _1420_ _2466_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9043__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8181_ _3358_ _3395_ _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5393_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7132_ _0732_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7249__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8446__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8446__B2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7063_ _1473_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7512__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6014_ _1375_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4483__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8749__A2 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5680__B2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7965_ _3200_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6916_ _1186_ _4092_ _2158_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7896_ _3139_ _4349_ _3140_ _3141_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_74_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6847_ _2128_ _2159_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_52_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _2063_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6932__A1 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ _1131_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8517_ _2693_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8448_ _3422_ _3652_ _3667_ _3271_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_124_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__A1 as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5499__B2 as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8379_ _1400_ _3499_ _3583_ _3601_ _0334_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6160__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8437__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6999__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5671__A1 _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5877__I _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__B2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__C _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7176__B2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9066__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__I _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7479__A2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_51_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8676__A1 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4956__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8428__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7100__A1 _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8872__B _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7403__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8600__A1 _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7750_ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4962_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6701_ _1987_ _1990_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7681_ _2931_ _2932_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4893_ _4259_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7167__A1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ as2650.r0\[2\] _1860_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _4118_ _1869_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6390__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8302_ _2782_ _3527_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ as2650.holding_reg\[3\] _0917_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8667__A1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6494_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8233_ _2789_ _3423_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4528__I0 as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5445_ _0849_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8419__A1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8164_ _1297_ _3356_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5376_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7115_ _1792_ _2392_ _2397_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8338__I _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8095_ _2586_ _2660_ _3325_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _2337_ _2338_ _4401_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7642__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8997_ _0108_ clknet_leaf_47_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _3187_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9089__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7158__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7879_ _0311_ _3123_ _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7845__C _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5708__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6905__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7953__I0 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4916__B1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7417__I _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8022__B _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__A1 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5365__C _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4519__I0 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__B1 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7330__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8926__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7881__A2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4695__A2 _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8248__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7152__I _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8830__A1 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6991__I _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7397__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7327__I _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8649__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7771__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5230_ _0599_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _0477_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7062__I _4448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A2 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8821__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5092_ as2650.r123\[3\]\[2\] _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8920_ _0031_ clknet_leaf_35_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8851_ _4001_ _0997_ _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_6__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7802_ _3050_ _3010_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5994_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5310__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5938__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8782_ _2993_ _1761_ _3937_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7733_ _2966_ _2983_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _4228_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8888__A1 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7664_ _2606_ _2888_ _2897_ _0306_ _2916_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4876_ _4283_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _1925_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7595_ net34 _2810_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7560__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8949__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7237__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6546_ _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6477_ as2650.stack\[6\]\[12\] _1790_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6115__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8216_ _3441_ _3442_ _3443_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5428_ as2650.r123\[0\]\[2\] _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7863__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8147_ _3358_ _3357_ _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ _0765_ _0766_ _4383_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8078_ _4367_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _1961_ _2323_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5220__I _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8879__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6986__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A1 _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9104__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7854__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A1 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8803__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8803__B2 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7610__I _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6290__A1 _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5130__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8031__A2 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7090__I0 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7766__B _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6593__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ _4269_ _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _4248_ _4251_ _4254_ _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6400_ _1479_ _1736_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7380_ _0417_ _2637_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ _4171_ _4180_ _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _4318_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8098__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9050_ _0147_ clknet_leaf_46_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6262_ _0933_ _1599_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7845__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8001_ _2352_ _1259_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5213_ _0608_ _0619_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _0877_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _0551_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A1 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5608__B2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8270__A2 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _0494_ _4419_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__A2 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8903_ _0014_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8022__A2 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8834_ _1346_ _3981_ _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8765_ as2650.stack\[4\]\[1\] _3926_ _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7781__A1 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__A2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5977_ _1300_ _1354_ _1359_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7781__B2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7716_ _1378_ _2898_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _4433_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8696_ _1794_ _3873_ _3879_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7647_ _2842_ _2804_ _2843_ _2841_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_100_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ _4448_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6336__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9127__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7578_ net35 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8089__A2 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _0662_ _1836_ _1843_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9179_ _0276_ clknet_leaf_69_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5215__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8261__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4822__A2 _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6575__A2 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A1 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7524__B2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__B1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5838__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8788__B1 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4964__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8252__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__A2 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4813__A2 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _0970_ _1298_ _1281_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _2191_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5831_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7763__A1 _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6566__A2 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5762_ _1062_ _1059_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8550_ _2693_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7501_ _1023_ _1035_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xclkbuf_leaf_6_wb_clk_i clknet_3_1__leaf_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4713_ _4293_ _4306_ _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7515__A1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8481_ _0700_ _3698_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5693_ _1090_ _0523_ _1097_ _0669_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7432_ _2648_ _2610_ _2688_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ as2650.ins_reg\[3\] _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7363_ as2650.pc\[0\] net7 _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4575_ as2650.ins_reg\[4\] _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9102_ _0199_ clknet_leaf_15_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6314_ _0475_ _1618_ _1652_ _1524_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7294_ _4411_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5829__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5829__B2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9033_ _0144_ clknet_leaf_9_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6245_ _1578_ _1427_ _1585_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8491__A2 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6176_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4501__B2 _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4874__I _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5127_ _4413_ _0526_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5057__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ _4386_ _0371_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8790__B _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A2 _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8817_ _0778_ _3959_ _3969_ _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7754__A1 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8081__I _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8748_ _3900_ _2177_ _3909_ as2650.r123\[2\]\[3\] _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8679_ _2295_ _3865_ _3868_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7809__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__A1 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4784__I _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_76_wb_clk_i clknet_3_0__leaf_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__B1 _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__I _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5548__C _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7763__C _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4959__I as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4731__A1 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ _1370_ _1404_ _1405_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6484__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8166__I _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8225__A2 _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7981_ _2497_ _2501_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7984__A1 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _1842_ _2241_ _2242_ _2099_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6863_ _2174_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7736__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8602_ net28 _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5814_ _4184_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6794_ _0896_ _1826_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8533_ _3748_ _3749_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5745_ _1121_ _0664_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8464_ _2782_ _3681_ _3682_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ _1079_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7415_ _0338_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4869__I _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4627_ _4057_ _4184_ _4188_ _4220_ _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_117_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8395_ _0395_ _3614_ _3616_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A1 _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7346_ _2594_ _2598_ _2604_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _4150_ _4077_ _4151_ _4070_ _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7277_ _2536_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4489_ _4082_ as2650.r123_2\[1\]\[6\] _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6475__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__A2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9016_ _0127_ clknet_leaf_30_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ _4357_ _4297_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A1 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5450__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A1 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6994__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput40 net40 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5269__A2 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__I _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6218__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7966__A1 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5441__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8391__A1 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7194__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8391__B2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _0916_ _0921_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8143__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8143__B2 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4689__I as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ _4148_ _4154_ _4176_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8982__CLK clknet_3_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8694__A2 _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7200_ as2650.stack\[2\]\[12\] _2462_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8180_ _3277_ _3397_ _3408_ _3170_ _3032_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5392_ _4208_ _0798_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7131_ _2408_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8446__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7062_ _4448_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6013_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5313__I _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8624__I _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7964_ _3199_ as2650.holding_reg\[7\] _3165_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _2184_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7895_ _3139_ _4428_ _2600_ _4432_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6144__I _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6846_ _4075_ _1865_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _2065_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8516_ _3688_ _0806_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5728_ _0523_ _0652_ _0808_ _0569_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_109_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4599__I _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8447_ _3663_ _3666_ _2816_ _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5659_ _1056_ _0840_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9107__D _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5499__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__I1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8378_ _3596_ _3600_ _3391_ _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ _1274_ net7 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8437__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6319__I _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A1 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8534__I _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__A1 _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7594__B _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8676__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__I1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_wb_clk_i clknet_3_3__leaf_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7100__A2 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A1 _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7939__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_7__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8600__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5414__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _4400_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6700_ _2011_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7680_ _2885_ _2889_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4892_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8364__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6631_ as2650.r0\[1\] _1857_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9010__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6562_ _0589_ _1865_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8301_ _3344_ _3502_ _3508_ _3258_ _3526_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5513_ _4206_ _0540_ _0919_ _0595_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5308__I _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _4293_ _0792_ _1809_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6678__A1 _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8232_ _1314_ _3272_ _3459_ _3161_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4528__I1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9160__CLK clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5444_ _0850_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8163_ _1298_ _3272_ _3392_ _3161_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5375_ net8 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7114_ as2650.stack\[4\]\[10\] _2395_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8094_ _2663_ _1692_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7045_ _4046_ _4270_ _1244_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5043__I _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8996_ _0107_ clknet_leaf_49_wb_clk_i as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7947_ _3185_ as2650.holding_reg\[3\] _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7878_ _4405_ _0345_ _2518_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8355__A1 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6829_ _1832_ _2111_ _2143_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8303__B _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7953__I1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4916__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__B2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__A2 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4519__I1 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__B2 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7330__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5341__A1 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7881__A3 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7618__B1 _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5381__C _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8830__A2 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6841__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4792__I _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8594__A1 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9033__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__A1 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__B2 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8897__A2 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6512__I _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9183__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4967__I _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5160_ _0523_ _0537_ _0544_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7085__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5091_ _0507_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8821__A2 _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6832__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8850_ _0925_ _0934_ _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7801_ net39 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8781_ _1680_ _1754_ _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5993_ _4360_ _0479_ _0560_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_64_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6060__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7732_ _2967_ _2953_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4944_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8337__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7663_ _2911_ _2912_ _2915_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4875_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8888__A2 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6899__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6422__I _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _1928_ _1930_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7594_ _2839_ _2847_ _0314_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7560__A2 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _4149_ _4159_ _1859_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5571__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5038__I _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6476_ _1419_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7312__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8215_ _2767_ _3396_ _2789_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5427_ _0747_ _0578_ _0835_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8146_ _3277_ _3360_ _3375_ _3032_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ _0765_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__B _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7076__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8077_ _1510_ _3308_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5289_ as2650.psu\[0\] _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__A1 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ _1909_ _1937_ _1960_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_102_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9056__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9120__D _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8576__A1 _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8979_ _0090_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8033__B _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8879__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7428__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7000__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__A3 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8500__A1 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8803__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8016__B1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5411__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__A1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7090__I1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8319__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6593__A3 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5567__B _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4660_ _4253_ _4226_ _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7542__A2 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5553__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _4095_ _4097_ _4101_ _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6330_ _1619_ _4156_ _1667_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6261_ _0922_ _0923_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7073__I _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8000_ _4050_ _3227_ _3231_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ _0607_ _0619_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1530_ _1543_ _1544_ _1508_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7058__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5143_ _4373_ _4319_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_111_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7801__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _4055_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8902_ _4043_ _4044_ _3648_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6281__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8558__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8833_ _1436_ _3983_ _3984_ _3939_ _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__A1 _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8916__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8764_ _2279_ _3925_ _3927_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5976_ as2650.stack\[1\]\[3\] _1355_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7781__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7715_ _1389_ _2840_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4927_ _0348_ _0349_ _0343_ _0352_ _0336_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_127_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8695_ as2650.stack\[5\]\[11\] _3876_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6152__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7646_ _2898_ _1154_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5196__C _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ _4450_ _4326_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6336__A3 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7692__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8730__B2 as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7577_ _2787_ _2828_ _2831_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__I _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4789_ _4382_ _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6528_ _1821_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6459_ _1348_ _1366_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5847__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9178_ _0275_ clknet_leaf_31_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__A1 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8129_ _2663_ _3335_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8797__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6272__A2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8549__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7524__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8721__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__I _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__B2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5406__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8788__A1 _4424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8788__B2 _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__A3 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__A2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__I _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7212__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _1231_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7763__A2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5761_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5774__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4577__A2 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7500_ _2650_ _2754_ _2689_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4712_ _4305_ _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8480_ _3697_ _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5692_ _1095_ _0788_ _1096_ _1026_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7431_ _0881_ _0874_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4643_ _4236_ _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8401__B _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7362_ _0324_ _2619_ _2599_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4574_ _4116_ _4126_ _4167_ _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9101_ _0198_ clknet_leaf_40_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7279__A1 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1122_ _0475_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7293_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9032_ _0143_ clknet_leaf_21_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6244_ as2650.stack\[3\]\[13\] _1576_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8491__A3 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _1517_ _1523_ _1526_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_58_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7531__I _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8779__A1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5126_ _0528_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7451__A1 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6147__I _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5057_ _4060_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_72_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__A1 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8816_ _3959_ _3968_ _0732_ _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8747_ _3915_ _3916_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5959_ _1331_ _1340_ _1345_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8678_ as2650.stack\[6\]\[5\] _3866_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8703__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7629_ _1320_ _1141_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4740__A2 _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8482__A3 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7690__A1 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7441__I _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7442__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6057__I as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__B2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_4__leaf_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6520__I _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7681__A1 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4975__I _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8891__B _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6236__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7980_ _4384_ _1266_ _2488_ _4327_ _3212_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7984__A2 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _4202_ _1842_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6862_ _2114_ _2140_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7736__A2 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8115__C _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8601_ _0815_ _3493_ _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5813_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5747__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6793_ _2097_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8532_ _1540_ _3731_ _2482_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5744_ _1028_ _0669_ _1147_ _0689_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8463_ _1429_ _1755_ _3670_ _3339_ _3555_ _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5675_ _4126_ _1011_ _4116_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7526__I _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7414_ _1588_ _2658_ _2662_ _4276_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6172__A1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _4198_ _4204_ _4219_ _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8394_ _3537_ _3604_ _3615_ _3235_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7970__B _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7345_ _4437_ _2599_ _2603_ _2549_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5046__I _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _4108_ _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4722__A2 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7276_ _1215_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4488_ _4063_ _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_85_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9015_ _0126_ clknet_leaf_35_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7672__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6475__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__A3 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4486__A1 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _4439_ _0445_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7424__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _4393_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6089_ as2650.r123_2\[3\]\[1\] _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A2 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6605__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7436__I _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__I _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6163__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput30 net30 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7663__A1 _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_3_3__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7966__A2 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6515__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5559__C _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8143__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6250__I _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _4191_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5391_ _0798_ _0654_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7130_ _2407_ _0815_ _1808_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7061_ _2353_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6012_ as2650.pc\[9\] _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

