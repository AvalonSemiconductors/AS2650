// This is the unpowered netlist.
module serial_ports (RXD,
    TXD,
    bus_cyc,
    bus_we,
    io_in,
    irq3,
    rst,
    wb_clk_i,
    addr,
    data_in,
    data_out,
    io_oeb,
    io_out);
 input RXD;
 output TXD;
 input bus_cyc;
 input bus_we;
 input io_in;
 output irq3;
 input rst;
 input wb_clk_i;
 input [2:0] addr;
 input [7:0] data_in;
 output [7:0] data_out;
 output [2:0] io_oeb;
 output [2:0] io_out;

 wire net29;
 wire net30;
 wire net32;
 wire net31;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \spi.busy ;
 wire \spi.counter[0] ;
 wire \spi.counter[1] ;
 wire \spi.counter[2] ;
 wire \spi.counter[3] ;
 wire \spi.counter[4] ;
 wire \spi.data_in_buff[0] ;
 wire \spi.data_in_buff[1] ;
 wire \spi.data_in_buff[2] ;
 wire \spi.data_in_buff[3] ;
 wire \spi.data_in_buff[4] ;
 wire \spi.data_in_buff[5] ;
 wire \spi.data_in_buff[6] ;
 wire \spi.data_in_buff[7] ;
 wire \spi.data_out_buff[0] ;
 wire \spi.data_out_buff[1] ;
 wire \spi.data_out_buff[2] ;
 wire \spi.data_out_buff[3] ;
 wire \spi.data_out_buff[4] ;
 wire \spi.data_out_buff[5] ;
 wire \spi.data_out_buff[6] ;
 wire \spi.data_out_buff[7] ;
 wire \spi.div_counter[0] ;
 wire \spi.div_counter[1] ;
 wire \spi.div_counter[2] ;
 wire \spi.div_counter[3] ;
 wire \spi.div_counter[4] ;
 wire \spi.div_counter[5] ;
 wire \spi.div_counter[6] ;
 wire \spi.div_counter[7] ;
 wire \spi.divisor[0] ;
 wire \spi.divisor[1] ;
 wire \spi.divisor[2] ;
 wire \spi.divisor[3] ;
 wire \spi.divisor[4] ;
 wire \spi.divisor[5] ;
 wire \spi.divisor[6] ;
 wire \spi.divisor[7] ;
 wire \spi.dout[0] ;
 wire \spi.dout[1] ;
 wire \spi.dout[2] ;
 wire \spi.dout[3] ;
 wire \spi.dout[4] ;
 wire \spi.dout[5] ;
 wire \spi.dout[6] ;
 wire \spi.dout[7] ;
 wire \uart.busy ;
 wire \uart.counter[0] ;
 wire \uart.counter[1] ;
 wire \uart.counter[2] ;
 wire \uart.counter[3] ;
 wire \uart.data_buff[0] ;
 wire \uart.data_buff[1] ;
 wire \uart.data_buff[2] ;
 wire \uart.data_buff[3] ;
 wire \uart.data_buff[4] ;
 wire \uart.data_buff[5] ;
 wire \uart.data_buff[6] ;
 wire \uart.data_buff[7] ;
 wire \uart.data_buff[8] ;
 wire \uart.data_buff[9] ;
 wire \uart.div_counter[0] ;
 wire \uart.div_counter[10] ;
 wire \uart.div_counter[11] ;
 wire \uart.div_counter[12] ;
 wire \uart.div_counter[13] ;
 wire \uart.div_counter[14] ;
 wire \uart.div_counter[15] ;
 wire \uart.div_counter[1] ;
 wire \uart.div_counter[2] ;
 wire \uart.div_counter[3] ;
 wire \uart.div_counter[4] ;
 wire \uart.div_counter[5] ;
 wire \uart.div_counter[6] ;
 wire \uart.div_counter[7] ;
 wire \uart.div_counter[8] ;
 wire \uart.div_counter[9] ;
 wire \uart.divisor[0] ;
 wire \uart.divisor[10] ;
 wire \uart.divisor[11] ;
 wire \uart.divisor[12] ;
 wire \uart.divisor[13] ;
 wire \uart.divisor[14] ;
 wire \uart.divisor[15] ;
 wire \uart.divisor[1] ;
 wire \uart.divisor[2] ;
 wire \uart.divisor[3] ;
 wire \uart.divisor[4] ;
 wire \uart.divisor[5] ;
 wire \uart.divisor[6] ;
 wire \uart.divisor[7] ;
 wire \uart.divisor[8] ;
 wire \uart.divisor[9] ;
 wire \uart.dout[0] ;
 wire \uart.dout[1] ;
 wire \uart.dout[2] ;
 wire \uart.dout[3] ;
 wire \uart.dout[4] ;
 wire \uart.dout[5] ;
 wire \uart.dout[6] ;
 wire \uart.dout[7] ;
 wire \uart.has_byte ;
 wire \uart.receive_buff[0] ;
 wire \uart.receive_buff[1] ;
 wire \uart.receive_buff[2] ;
 wire \uart.receive_buff[3] ;
 wire \uart.receive_buff[4] ;
 wire \uart.receive_buff[5] ;
 wire \uart.receive_buff[6] ;
 wire \uart.receive_buff[7] ;
 wire \uart.receive_counter[0] ;
 wire \uart.receive_counter[1] ;
 wire \uart.receive_counter[2] ;
 wire \uart.receive_counter[3] ;
 wire \uart.receive_div_counter[0] ;
 wire \uart.receive_div_counter[10] ;
 wire \uart.receive_div_counter[11] ;
 wire \uart.receive_div_counter[12] ;
 wire \uart.receive_div_counter[13] ;
 wire \uart.receive_div_counter[14] ;
 wire \uart.receive_div_counter[15] ;
 wire \uart.receive_div_counter[1] ;
 wire \uart.receive_div_counter[2] ;
 wire \uart.receive_div_counter[3] ;
 wire \uart.receive_div_counter[4] ;
 wire \uart.receive_div_counter[5] ;
 wire \uart.receive_div_counter[6] ;
 wire \uart.receive_div_counter[7] ;
 wire \uart.receive_div_counter[8] ;
 wire \uart.receive_div_counter[9] ;
 wire \uart.receiving ;
 wire uart_ien;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__I (.I(\spi.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0834__I (.I(\spi.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0836__A1 (.I(\spi.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0836__B2 (.I(\spi.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0840__A1 (.I(\spi.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0842__A1 (.I(\spi.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0842__B2 (.I(\spi.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0846__A1 (.I(\spi.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0854__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0855__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0857__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0858__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0858__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0860__I (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0862__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0863__I (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0864__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0866__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0867__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0870__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0875__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0881__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0888__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0901__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0905__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0906__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__A1 (.I(\spi.data_out_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0915__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0919__A3 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0944__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0948__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0951__I (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0954__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__C (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0968__B (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0972__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0973__C (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0982__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0987__B (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__B (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__B (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__B (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A2 (.I(\spi.data_out_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1007__C (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__B (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1015__B (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1016__I (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1033__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1035__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1037__I0 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1039__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1039__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1040__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1041__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1045__A1 (.I(\uart.divisor[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1046__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1047__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1048__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1049__A1 (.I(\uart.divisor[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1051__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1055__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1056__A1 (.I(\uart.divisor[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1060__A1 (.I(\uart.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1062__I (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1064__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1066__A1 (.I(\uart.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1069__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1070__A1 (.I(\uart.divisor[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1073__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1074__A1 (.I(\uart.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1077__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1078__A1 (.I(\uart.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__A3 (.I(\uart.has_byte ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1081__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1085__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1088__A1 (.I(\uart.divisor[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1089__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1091__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1092__B1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1092__B2 (.I(\uart.divisor[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1095__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1097__I (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1098__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1100__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1102__B2 (.I(\uart.busy ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1103__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1105__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1107__A1 (.I(\uart.divisor[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1107__B1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1107__B2 (.I(\uart.divisor[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1111__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1113__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1114__B (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1115__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1116__A1 (.I(\uart.divisor[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1116__B1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1116__B2 (.I(\uart.divisor[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1118__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1119__B2 (.I(\uart.has_byte ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1120__B (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1121__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1124__I (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1125__B1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1126__A1 (.I(\uart.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1126__B2 (.I(\spi.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1129__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1131__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1134__A1 (.I(\uart.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1134__B2 (.I(\spi.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1135__A3 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1137__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1138__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1139__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1142__A1 (.I(\uart.divisor[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1143__A3 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1148__A1 (.I(\uart.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1148__B2 (.I(\spi.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1149__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1149__A3 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1153__B2 (.I(\uart.divisor[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1154__A1 (.I(\uart.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1154__B2 (.I(\spi.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1155__A1 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1155__A3 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1160__A2 (.I(\uart.divisor[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__A2 (.I(\uart.divisor[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__A2 (.I(\uart.divisor[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1167__A2 (.I(\uart.divisor[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__A2 (.I(\uart.divisor[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1171__A2 (.I(\uart.divisor[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__A2 (.I(\uart.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1173__A2 (.I(\uart.divisor[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__A1 (.I(\uart.receive_div_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1175__A2 (.I(\uart.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1176__A2 (.I(\uart.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1177__A2 (.I(\uart.divisor[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__A2 (.I(\uart.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1181__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1187__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1192__A3 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1193__B (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1198__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1200__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1202__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1205__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__A1 (.I(\uart.divisor[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1210__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1210__C (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__A1 (.I(\uart.divisor[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1212__C (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1214__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__A1 (.I(\uart.divisor[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1217__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1218__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1220__B (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1222__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1229__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1233__A1 (.I(\uart.divisor[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1244__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1249__A1 (.I(\spi.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1251__B (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1254__B (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__B (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1258__A1 (.I(\spi.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__B (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1263__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1264__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1267__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1278__B (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1280__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1293__C (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1296__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1297__B (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1299__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1308__B (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1313__A1 (.I(\uart.receive_div_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1314__I (.I(\uart.receive_div_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1317__A1 (.I(\uart.receive_div_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1322__B (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1333__B (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1337__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1342__B (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1345__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1347__B (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__B (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1357__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__B (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__B (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1387__B (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1389__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A1 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__A2 (.I(\uart.divisor[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1395__A2 (.I(\uart.divisor[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__A2 (.I(\uart.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A1 (.I(\uart.div_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A2 (.I(\uart.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1401__A2 (.I(\uart.divisor[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A2 (.I(\uart.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1406__A2 (.I(\uart.divisor[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A2 (.I(\uart.divisor[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A2 (.I(\uart.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A1 (.I(\uart.div_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__A2 (.I(\uart.divisor[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1413__A2 (.I(\uart.divisor[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1414__A2 (.I(\uart.divisor[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1419__A1 (.I(\uart.busy ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1421__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1427__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1429__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__C (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__I (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__B (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__C (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__B (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1460__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1460__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1466__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__C (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1491__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A1 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__B (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__B (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__B (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__I (.I(\uart.div_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A1 (.I(\uart.div_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A1 (.I(\uart.div_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A1 (.I(\uart.div_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__C (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A1 (.I(\uart.has_byte ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__B (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__C (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A2 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A2 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A2 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1663__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1671__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__CLK (.I(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__CLK (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__CLK (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__CLK (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__CLK (.I(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__CLK (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__CLK (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__CLK (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__CLK (.I(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__CLK (.I(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__CLK (.I(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__CLK (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__CLK (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__CLK (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__CLK (.I(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__CLK (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__CLK (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__CLK (.I(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__CLK (.I(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__CLK (.I(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__CLK (.I(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__CLK (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__D (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1782__CLK (.I(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__CLK (.I(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__CLK (.I(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__CLK (.I(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(RXD));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0827_ (.I(net16),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0828_ (.I(_0244_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0829_ (.I(_0245_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0830_ (.I(\spi.counter[0] ),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0831_ (.I(\spi.div_counter[7] ),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0832_ (.I(\spi.div_counter[4] ),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0833_ (.I(\spi.divisor[6] ),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0834_ (.I(\spi.divisor[3] ),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0835_ (.A1(_0250_),
    .A2(\spi.div_counter[6] ),
    .B1(\spi.div_counter[3] ),
    .B2(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _0836_ (.A1(\spi.divisor[7] ),
    .A2(_0248_),
    .B1(_0249_),
    .B2(\spi.divisor[4] ),
    .C(_0252_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0837_ (.I(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0838_ (.I(\spi.div_counter[2] ),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0839_ (.I(\spi.divisor[2] ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0840_ (.A1(\spi.divisor[7] ),
    .A2(_0248_),
    .B1(_0255_),
    .B2(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0841_ (.I(\spi.div_counter[6] ),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0842_ (.A1(\spi.divisor[6] ),
    .A2(_0258_),
    .B1(_0249_),
    .B2(\spi.divisor[4] ),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0843_ (.I(\spi.div_counter[3] ),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0844_ (.I(\spi.div_counter[2] ),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0845_ (.A1(\spi.divisor[0] ),
    .A2(\spi.div_counter[0] ),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0846_ (.A1(\spi.divisor[3] ),
    .A2(_0260_),
    .B1(_0261_),
    .B2(\spi.divisor[2] ),
    .C(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0847_ (.A1(\spi.divisor[1] ),
    .A2(\spi.div_counter[1] ),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0848_ (.A1(\spi.divisor[5] ),
    .A2(\spi.div_counter[5] ),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0849_ (.A1(_0264_),
    .A2(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0850_ (.A1(_0257_),
    .A2(_0259_),
    .A3(_0263_),
    .A4(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0851_ (.I(_0267_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0852_ (.A1(_0247_),
    .A2(_0254_),
    .A3(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0853_ (.I(_0269_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0854_ (.I(net4),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0855_ (.I(net3),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0856_ (.I(_0272_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0857_ (.A1(_0273_),
    .A2(net2),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0858_ (.A1(net5),
    .A2(net6),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0859_ (.A1(_0271_),
    .A2(\spi.busy ),
    .A3(_0274_),
    .A4(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0860_ (.I(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0861_ (.I(_0277_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0862_ (.I(net7),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0863_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0864_ (.A1(_0280_),
    .A2(_0278_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0865_ (.A1(\spi.data_out_buff[0] ),
    .A2(_0278_),
    .B(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0866_ (.A1(_0246_),
    .A2(_0270_),
    .A3(_0282_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0867_ (.I(net16),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0868_ (.I(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0869_ (.I(_0284_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0870_ (.I(net8),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0871_ (.I(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0872_ (.I(_0277_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0873_ (.A1(\spi.data_out_buff[1] ),
    .A2(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0874_ (.I(_0269_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0875_ (.A1(_0287_),
    .A2(_0278_),
    .B(_0289_),
    .C(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0876_ (.A1(\spi.data_out_buff[0] ),
    .A2(_0270_),
    .B(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0877_ (.A1(_0285_),
    .A2(_0292_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0878_ (.I(_0271_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0879_ (.A1(_0293_),
    .A2(\spi.busy ),
    .A3(_0274_),
    .A4(_0275_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0880_ (.I(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0881_ (.A1(\spi.data_out_buff[2] ),
    .A2(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0882_ (.I(_0277_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0883_ (.A1(net9),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0884_ (.I(_0269_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0885_ (.A1(_0296_),
    .A2(_0298_),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0886_ (.A1(\spi.data_out_buff[1] ),
    .A2(_0270_),
    .B(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0887_ (.A1(_0285_),
    .A2(_0301_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0888_ (.A1(\spi.data_out_buff[3] ),
    .A2(_0295_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0889_ (.A1(net10),
    .A2(_0297_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0890_ (.A1(_0302_),
    .A2(_0303_),
    .B(_0299_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0891_ (.A1(\spi.data_out_buff[2] ),
    .A2(_0270_),
    .B(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0892_ (.A1(_0285_),
    .A2(_0305_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0893_ (.I(_0269_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0894_ (.A1(\spi.data_out_buff[4] ),
    .A2(_0295_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0895_ (.A1(net11),
    .A2(_0297_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0896_ (.A1(_0307_),
    .A2(_0308_),
    .B(_0299_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0897_ (.A1(\spi.data_out_buff[3] ),
    .A2(_0306_),
    .B(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0898_ (.A1(_0285_),
    .A2(_0310_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0899_ (.I(_0284_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0900_ (.I(_0294_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0901_ (.A1(\spi.data_out_buff[5] ),
    .A2(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0902_ (.A1(net12),
    .A2(_0288_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0903_ (.A1(_0313_),
    .A2(_0314_),
    .B(_0290_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0904_ (.A1(\spi.data_out_buff[4] ),
    .A2(_0306_),
    .B(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0905_ (.A1(_0311_),
    .A2(_0316_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0906_ (.A1(\spi.data_out_buff[6] ),
    .A2(_0312_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0907_ (.A1(net13),
    .A2(_0288_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0908_ (.A1(_0317_),
    .A2(_0318_),
    .B(_0290_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0909_ (.A1(\spi.data_out_buff[5] ),
    .A2(_0306_),
    .B(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0910_ (.A1(_0311_),
    .A2(_0320_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0911_ (.A1(\spi.data_out_buff[7] ),
    .A2(_0312_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0912_ (.A1(net14),
    .A2(_0288_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0913_ (.A1(_0321_),
    .A2(_0322_),
    .B(_0290_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0914_ (.A1(\spi.data_out_buff[6] ),
    .A2(_0306_),
    .B(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0915_ (.A1(_0311_),
    .A2(_0324_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0916_ (.A1(\spi.counter[0] ),
    .A2(\spi.counter[1] ),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0917_ (.A1(\spi.counter[2] ),
    .A2(\spi.counter[3] ),
    .A3(\spi.counter[4] ),
    .A4(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0918_ (.I(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0919_ (.A1(_0254_),
    .A2(_0268_),
    .A3(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0920_ (.A1(_0297_),
    .A2(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0921_ (.I(_0283_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0922_ (.A1(_0247_),
    .A2(_0329_),
    .B(_0299_),
    .C(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0923_ (.I(_0331_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0924_ (.I(\spi.counter[1] ),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0925_ (.I(\spi.counter[0] ),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0926_ (.A1(_0333_),
    .A2(_0332_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0927_ (.I(_0328_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0928_ (.A1(_0332_),
    .A2(_0329_),
    .B1(_0334_),
    .B2(_0335_),
    .C(_0330_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0929_ (.I(_0336_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0930_ (.I(\spi.counter[2] ),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0931_ (.A1(_0247_),
    .A2(_0332_),
    .A3(_0337_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0932_ (.A1(_0247_),
    .A2(_0332_),
    .B(_0337_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0933_ (.A1(_0338_),
    .A2(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0934_ (.A1(_0337_),
    .A2(_0329_),
    .B1(_0340_),
    .B2(_0335_),
    .C(_0330_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0935_ (.I(_0341_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0936_ (.I(\spi.counter[3] ),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0937_ (.A1(_0342_),
    .A2(_0338_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0938_ (.A1(_0342_),
    .A2(_0329_),
    .B1(_0343_),
    .B2(_0335_),
    .C(_0330_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0939_ (.I(_0344_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0940_ (.I(_0244_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0941_ (.I(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0942_ (.A1(_0254_),
    .A2(_0268_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0943_ (.A1(_0337_),
    .A2(\spi.counter[3] ),
    .A3(\spi.counter[4] ),
    .A4(_0325_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0944_ (.A1(_0347_),
    .A2(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0945_ (.A1(_0342_),
    .A2(\spi.counter[4] ),
    .A3(_0349_),
    .A4(_0338_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0946_ (.A1(_0342_),
    .A2(_0349_),
    .A3(_0338_),
    .B(\spi.counter[4] ),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0947_ (.A1(_0254_),
    .A2(_0268_),
    .B(_0278_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0948_ (.A1(_0346_),
    .A2(_0350_),
    .A3(_0351_),
    .A4(_0352_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0949_ (.I(_0244_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0950_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0951_ (.I(_0327_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0952_ (.I(_0355_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0953_ (.I(_0283_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0954_ (.A1(\spi.busy ),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0955_ (.A1(_0354_),
    .A2(_0356_),
    .B(_0358_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0956_ (.I(\spi.div_counter[0] ),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0957_ (.A1(_0312_),
    .A2(_0327_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0958_ (.A1(_0347_),
    .A2(_0326_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0959_ (.I(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0960_ (.A1(_0359_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0961_ (.A1(_0359_),
    .A2(_0360_),
    .B(_0363_),
    .C(_0354_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0962_ (.I(\spi.div_counter[1] ),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0963_ (.A1(_0277_),
    .A2(_0348_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0964_ (.I(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0965_ (.A1(_0364_),
    .A2(_0359_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0966_ (.A1(_0364_),
    .A2(_0366_),
    .B1(_0362_),
    .B2(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0967_ (.I(_0345_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0968_ (.A1(_0364_),
    .A2(_0359_),
    .B(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0969_ (.A1(_0368_),
    .A2(_0370_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0970_ (.A1(_0255_),
    .A2(_0364_),
    .A3(\spi.div_counter[0] ),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0971_ (.A1(_0255_),
    .A2(_0365_),
    .B1(_0361_),
    .B2(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0972_ (.I(_0353_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0973_ (.A1(_0261_),
    .A2(_0367_),
    .B(_0372_),
    .C(_0373_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0974_ (.I(_0361_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0975_ (.A1(_0260_),
    .A2(_0371_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0976_ (.A1(\spi.div_counter[3] ),
    .A2(_0366_),
    .B1(_0374_),
    .B2(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0977_ (.A1(_0311_),
    .A2(_0376_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0978_ (.I(_0284_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0979_ (.A1(\spi.div_counter[3] ),
    .A2(_0255_),
    .A3(\spi.div_counter[1] ),
    .A4(\spi.div_counter[0] ),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0980_ (.A1(\spi.div_counter[4] ),
    .A2(_0378_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0981_ (.A1(\spi.div_counter[4] ),
    .A2(_0366_),
    .B1(_0374_),
    .B2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0982_ (.A1(_0377_),
    .A2(_0380_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0983_ (.I(\spi.div_counter[5] ),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0984_ (.A1(\spi.div_counter[4] ),
    .A2(_0378_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0985_ (.A1(_0381_),
    .A2(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0986_ (.A1(_0381_),
    .A2(_0366_),
    .B1(_0362_),
    .B2(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0987_ (.A1(_0381_),
    .A2(_0382_),
    .B(_0369_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0988_ (.A1(_0384_),
    .A2(_0385_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0989_ (.A1(_0258_),
    .A2(_0381_),
    .A3(_0362_),
    .A4(_0382_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0990_ (.A1(_0258_),
    .A2(_0383_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0991_ (.A1(_0347_),
    .A2(_0355_),
    .A3(_0387_),
    .B(_0360_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0992_ (.A1(\spi.div_counter[6] ),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0993_ (.I(_0244_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0994_ (.I(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0995_ (.A1(_0386_),
    .A2(_0389_),
    .B(_0391_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0996_ (.A1(\spi.div_counter[7] ),
    .A2(_0388_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0997_ (.A1(_0248_),
    .A2(_0374_),
    .A3(_0387_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0998_ (.A1(_0392_),
    .A2(_0393_),
    .B(_0391_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0999_ (.A1(_0333_),
    .A2(_0253_),
    .A3(_0267_),
    .A4(_0326_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1000_ (.I(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1001_ (.I(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1002_ (.A1(_0284_),
    .A2(_0374_),
    .A3(_0396_),
    .B(net27),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1003_ (.A1(_0333_),
    .A2(\spi.data_out_buff[7] ),
    .A3(_0369_),
    .A4(_0335_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1004_ (.A1(_0397_),
    .A2(_0398_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1005_ (.I(\spi.data_in_buff[0] ),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1006_ (.A1(\spi.dout[0] ),
    .A2(_0355_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1007_ (.A1(_0399_),
    .A2(_0356_),
    .B(_0400_),
    .C(_0373_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1008_ (.A1(\spi.data_in_buff[1] ),
    .A2(_0356_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1009_ (.I(_0348_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1010_ (.I(_0402_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1011_ (.A1(\spi.dout[1] ),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1012_ (.A1(_0401_),
    .A2(_0404_),
    .B(_0391_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1013_ (.A1(\spi.data_in_buff[2] ),
    .A2(_0356_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1014_ (.A1(\spi.dout[2] ),
    .A2(_0403_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1015_ (.A1(_0405_),
    .A2(_0406_),
    .B(_0391_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1016_ (.I(_0327_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1017_ (.A1(\spi.data_in_buff[3] ),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1018_ (.A1(\spi.dout[3] ),
    .A2(_0403_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1019_ (.I(_0390_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1020_ (.A1(_0408_),
    .A2(_0409_),
    .B(_0410_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1021_ (.A1(\spi.data_in_buff[4] ),
    .A2(_0407_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1022_ (.A1(\spi.dout[4] ),
    .A2(_0403_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1023_ (.A1(_0411_),
    .A2(_0412_),
    .B(_0410_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1024_ (.A1(\spi.data_in_buff[5] ),
    .A2(_0407_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1025_ (.A1(\spi.dout[5] ),
    .A2(_0402_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1026_ (.A1(_0413_),
    .A2(_0414_),
    .B(_0410_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1027_ (.A1(\spi.data_in_buff[6] ),
    .A2(_0407_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1028_ (.A1(\spi.dout[6] ),
    .A2(_0402_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1029_ (.A1(_0415_),
    .A2(_0416_),
    .B(_0410_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1030_ (.A1(\spi.data_in_buff[7] ),
    .A2(_0355_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1031_ (.A1(\spi.dout[7] ),
    .A2(_0402_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1032_ (.I(net16),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1033_ (.I(_0419_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1034_ (.I(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1035_ (.A1(_0417_),
    .A2(_0418_),
    .B(_0421_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1036_ (.A1(_0295_),
    .A2(_0361_),
    .B(_0283_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1037_ (.I0(net26),
    .I1(_0396_),
    .S(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1038_ (.I(_0423_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1039_ (.A1(net5),
    .A2(net6),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1040_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1041_ (.I(net4),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1042_ (.A1(_0426_),
    .A2(_0274_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1043_ (.A1(_0425_),
    .A2(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1044_ (.I(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1045_ (.A1(\uart.divisor[0] ),
    .A2(_0428_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1046_ (.I(_0345_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1047_ (.I(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1048_ (.A1(_0280_),
    .A2(_0429_),
    .B(_0430_),
    .C(_0432_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1049_ (.A1(\uart.divisor[1] ),
    .A2(_0428_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1050_ (.A1(_0287_),
    .A2(_0429_),
    .B(_0433_),
    .C(_0432_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1051_ (.I(_0431_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1052_ (.I(net9),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1053_ (.A1(_0426_),
    .A2(_0274_),
    .A3(_0275_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1054_ (.I(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1055_ (.A1(_0435_),
    .A2(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1056_ (.A1(\uart.divisor[2] ),
    .A2(_0429_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1057_ (.A1(_0434_),
    .A2(_0438_),
    .A3(_0439_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1058_ (.I(net10),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1059_ (.A1(_0440_),
    .A2(_0437_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1060_ (.A1(\uart.divisor[3] ),
    .A2(_0429_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1061_ (.A1(_0434_),
    .A2(_0441_),
    .A3(_0442_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1062_ (.I(_0431_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1063_ (.I(net11),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1064_ (.A1(_0444_),
    .A2(_0437_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1065_ (.I(_0428_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1066_ (.A1(\uart.divisor[4] ),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1067_ (.A1(_0443_),
    .A2(_0445_),
    .A3(_0447_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1068_ (.I(net12),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1069_ (.A1(_0448_),
    .A2(_0437_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1070_ (.A1(\uart.divisor[5] ),
    .A2(_0446_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1071_ (.A1(_0443_),
    .A2(_0449_),
    .A3(_0450_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1072_ (.I(net13),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1073_ (.A1(_0451_),
    .A2(_0436_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1074_ (.A1(\uart.divisor[6] ),
    .A2(_0446_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1075_ (.A1(_0443_),
    .A2(_0452_),
    .A3(_0453_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1076_ (.I(net14),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1077_ (.A1(_0454_),
    .A2(_0436_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1078_ (.A1(\uart.divisor[7] ),
    .A2(_0446_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1079_ (.A1(_0443_),
    .A2(_0455_),
    .A3(_0456_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1080_ (.A1(uart_ien),
    .A2(_0346_),
    .A3(\uart.has_byte ),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1081_ (.I(_0457_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1082_ (.I(net5),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1083_ (.I(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1084_ (.I(_0427_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1085_ (.I(net2),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1086_ (.A1(_0293_),
    .A2(_0273_),
    .A3(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1087_ (.I(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1088_ (.A1(\uart.divisor[0] ),
    .A2(_0460_),
    .B1(_0463_),
    .B2(\uart.dout[0] ),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1089_ (.A1(_0426_),
    .A2(net3),
    .A3(_0461_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1090_ (.A1(_0426_),
    .A2(_0273_),
    .A3(_0461_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1091_ (.I(_0466_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1092_ (.A1(uart_ien),
    .A2(_0465_),
    .B1(_0467_),
    .B2(\uart.divisor[8] ),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1093_ (.A1(_0464_),
    .A2(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1094_ (.I(_0458_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1095_ (.I(net2),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1096_ (.A1(_0293_),
    .A2(_0273_),
    .A3(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1097_ (.I(_0472_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1098_ (.A1(net4),
    .A2(_0272_),
    .A3(_0471_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _1099_ (.I(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1100_ (.A1(_0293_),
    .A2(net3),
    .A3(_0461_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1101_ (.I(_0476_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1102_ (.A1(\spi.dout[0] ),
    .A2(_0473_),
    .B1(_0475_),
    .B2(\uart.busy ),
    .C1(_0477_),
    .C2(\spi.divisor[0] ),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1103_ (.A1(_0470_),
    .A2(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1104_ (.A1(_0459_),
    .A2(net18),
    .B1(_0469_),
    .B2(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1105_ (.A1(_0377_),
    .A2(_0480_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1106_ (.I(_0462_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _1107_ (.A1(\uart.divisor[1] ),
    .A2(_0460_),
    .B1(_0467_),
    .B2(\uart.divisor[9] ),
    .C1(\uart.dout[1] ),
    .C2(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1108_ (.I(_0476_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1109_ (.I(_0458_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1110_ (.A1(\spi.dout[1] ),
    .A2(_0473_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1111_ (.A1(_0484_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1112_ (.A1(\spi.divisor[1] ),
    .A2(_0483_),
    .B1(_0475_),
    .B2(\spi.busy ),
    .C(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1113_ (.I(_0345_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1114_ (.A1(_0459_),
    .A2(net19),
    .B(_0488_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1115_ (.A1(_0482_),
    .A2(_0487_),
    .B(_0489_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _1116_ (.A1(\uart.divisor[2] ),
    .A2(_0460_),
    .B1(_0467_),
    .B2(\uart.divisor[10] ),
    .C1(\uart.dout[2] ),
    .C2(_0481_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1117_ (.A1(\spi.dout[2] ),
    .A2(_0473_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1118_ (.A1(_0484_),
    .A2(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1119_ (.A1(\spi.divisor[2] ),
    .A2(_0483_),
    .B1(_0475_),
    .B2(\uart.has_byte ),
    .C(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1120_ (.A1(_0459_),
    .A2(net20),
    .B(_0488_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1121_ (.A1(_0490_),
    .A2(_0493_),
    .B(_0494_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1122_ (.I(_0458_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1123_ (.A1(\uart.dout[3] ),
    .A2(_0481_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1124_ (.I(_0472_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1125_ (.A1(\spi.dout[3] ),
    .A2(_0497_),
    .B1(_0467_),
    .B2(\uart.divisor[11] ),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1126_ (.A1(\uart.divisor[3] ),
    .A2(_0460_),
    .B1(_0483_),
    .B2(\spi.divisor[3] ),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1127_ (.A1(_0470_),
    .A2(_0496_),
    .A3(_0498_),
    .A4(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1128_ (.A1(_0495_),
    .A2(net21),
    .B(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1129_ (.A1(_0377_),
    .A2(_0501_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1130_ (.A1(\uart.dout[4] ),
    .A2(_0481_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1131_ (.I(_0466_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1132_ (.A1(\spi.dout[4] ),
    .A2(_0497_),
    .B1(_0503_),
    .B2(\uart.divisor[12] ),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1133_ (.I(_0427_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1134_ (.A1(\uart.divisor[4] ),
    .A2(_0505_),
    .B1(_0483_),
    .B2(\spi.divisor[4] ),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1135_ (.A1(_0470_),
    .A2(_0502_),
    .A3(_0504_),
    .A4(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1136_ (.A1(_0495_),
    .A2(net22),
    .B(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1137_ (.A1(_0377_),
    .A2(_0508_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1138_ (.I(_0419_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1139_ (.I(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1140_ (.A1(\uart.dout[5] ),
    .A2(_0463_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1141_ (.A1(\spi.dout[5] ),
    .A2(_0497_),
    .B1(_0503_),
    .B2(\uart.divisor[13] ),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1142_ (.A1(\uart.divisor[5] ),
    .A2(_0505_),
    .B1(_0477_),
    .B2(\spi.divisor[5] ),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1143_ (.A1(_0470_),
    .A2(_0511_),
    .A3(_0512_),
    .A4(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1144_ (.A1(_0495_),
    .A2(net23),
    .B(_0514_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1145_ (.A1(_0510_),
    .A2(_0515_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1146_ (.A1(\uart.dout[6] ),
    .A2(_0463_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1147_ (.A1(\spi.dout[6] ),
    .A2(_0497_),
    .B1(_0503_),
    .B2(\uart.divisor[14] ),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1148_ (.A1(\uart.divisor[6] ),
    .A2(_0505_),
    .B1(_0477_),
    .B2(\spi.divisor[6] ),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1149_ (.A1(_0484_),
    .A2(_0516_),
    .A3(_0517_),
    .A4(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1150_ (.A1(_0459_),
    .A2(net24),
    .B(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1151_ (.A1(_0510_),
    .A2(_0520_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1152_ (.A1(\uart.dout[7] ),
    .A2(_0463_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1153_ (.A1(\spi.dout[7] ),
    .A2(_0473_),
    .B1(_0503_),
    .B2(\uart.divisor[15] ),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1154_ (.A1(\uart.divisor[7] ),
    .A2(_0505_),
    .B1(_0477_),
    .B2(\spi.divisor[7] ),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1155_ (.A1(_0484_),
    .A2(_0521_),
    .A3(_0522_),
    .A4(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1156_ (.A1(net25),
    .A2(_0495_),
    .B(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1157_ (.A1(_0510_),
    .A2(_0525_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1158_ (.I(\uart.receiving ),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1159_ (.A1(\uart.receive_div_counter[14] ),
    .A2(\uart.divisor[14] ),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1160_ (.A1(\uart.receive_div_counter[9] ),
    .A2(\uart.divisor[9] ),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1161_ (.A1(\uart.receive_div_counter[12] ),
    .A2(\uart.divisor[12] ),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1162_ (.A1(\uart.receive_div_counter[10] ),
    .A2(\uart.divisor[10] ),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1163_ (.A1(_0527_),
    .A2(_0528_),
    .A3(_0529_),
    .A4(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1164_ (.A1(\uart.receive_div_counter[13] ),
    .A2(\uart.divisor[13] ),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1165_ (.A1(\uart.receive_div_counter[1] ),
    .A2(\uart.divisor[1] ),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1166_ (.A1(\uart.receive_div_counter[11] ),
    .A2(\uart.divisor[11] ),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1167_ (.A1(\uart.receive_div_counter[15] ),
    .A2(\uart.divisor[15] ),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1168_ (.A1(_0532_),
    .A2(_0533_),
    .A3(_0534_),
    .A4(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1169_ (.A1(_0531_),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1170_ (.A1(\uart.receive_div_counter[0] ),
    .A2(\uart.divisor[0] ),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1171_ (.A1(\uart.receive_div_counter[8] ),
    .A2(\uart.divisor[8] ),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1172_ (.A1(\uart.receive_div_counter[6] ),
    .A2(\uart.divisor[6] ),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1173_ (.A1(\uart.receive_div_counter[5] ),
    .A2(\uart.divisor[5] ),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1174_ (.A1(_0538_),
    .A2(_0539_),
    .A3(_0540_),
    .A4(_0541_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1175_ (.A1(\uart.receive_div_counter[7] ),
    .A2(\uart.divisor[7] ),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1176_ (.A1(\uart.receive_div_counter[4] ),
    .A2(\uart.divisor[4] ),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1177_ (.A1(\uart.receive_div_counter[2] ),
    .A2(\uart.divisor[2] ),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1178_ (.A1(\uart.receive_div_counter[3] ),
    .A2(\uart.divisor[3] ),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1179_ (.A1(_0543_),
    .A2(_0544_),
    .A3(_0545_),
    .A4(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1180_ (.A1(_0542_),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1181_ (.A1(_0526_),
    .A2(_0537_),
    .A3(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1182_ (.A1(\uart.receive_counter[0] ),
    .A2(_0549_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1183_ (.I(_0526_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1184_ (.I(net1),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1185_ (.A1(_0551_),
    .A2(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1186_ (.A1(\uart.receive_counter[0] ),
    .A2(_0549_),
    .A3(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1187_ (.A1(_0550_),
    .A2(_0554_),
    .B(_0421_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1188_ (.A1(\uart.receive_counter[1] ),
    .A2(_0553_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1189_ (.A1(_0550_),
    .A2(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1190_ (.A1(_0510_),
    .A2(_0556_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1191_ (.A1(\uart.receive_counter[2] ),
    .A2(_0553_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1192_ (.A1(\uart.receive_counter[1] ),
    .A2(\uart.receive_counter[0] ),
    .A3(_0549_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1193_ (.A1(_0557_),
    .A2(_0558_),
    .B(_0488_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1194_ (.A1(_0557_),
    .A2(_0558_),
    .B(_0559_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1195_ (.I(\uart.receive_counter[3] ),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1196_ (.A1(_0560_),
    .A2(_0553_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1197_ (.A1(\uart.receive_counter[1] ),
    .A2(\uart.receive_counter[0] ),
    .A3(\uart.receive_counter[2] ),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1198_ (.A1(_0549_),
    .A2(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1199_ (.A1(_0561_),
    .A2(_0563_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1200_ (.A1(_0346_),
    .A2(_0564_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1201_ (.I(_0565_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1202_ (.A1(_0424_),
    .A2(_0465_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1203_ (.A1(_0286_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1204_ (.I0(net7),
    .I1(uart_ien),
    .S(_0567_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1205_ (.A1(_0346_),
    .A2(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1206_ (.I(_0569_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1207_ (.A1(_0424_),
    .A2(_0466_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1208_ (.I(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1209_ (.A1(\uart.divisor[8] ),
    .A2(_0570_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1210_ (.A1(_0280_),
    .A2(_0571_),
    .B(_0572_),
    .C(_0373_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1211_ (.A1(\uart.divisor[9] ),
    .A2(_0570_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1212_ (.A1(_0287_),
    .A2(_0571_),
    .B(_0573_),
    .C(_0373_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1213_ (.A1(_0435_),
    .A2(_0571_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1214_ (.A1(_0425_),
    .A2(_0466_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1215_ (.I(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1216_ (.A1(\uart.divisor[10] ),
    .A2(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1217_ (.A1(_0574_),
    .A2(_0577_),
    .B(_0421_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1218_ (.A1(_0440_),
    .A2(_0571_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1219_ (.A1(\uart.divisor[11] ),
    .A2(_0576_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1220_ (.A1(_0578_),
    .A2(_0579_),
    .B(_0421_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1221_ (.I(_0570_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1222_ (.A1(_0444_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1223_ (.A1(\uart.divisor[12] ),
    .A2(_0576_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1224_ (.I(_0420_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1225_ (.A1(_0581_),
    .A2(_0582_),
    .B(_0583_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1226_ (.A1(_0448_),
    .A2(_0580_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1227_ (.A1(\uart.divisor[13] ),
    .A2(_0576_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1228_ (.A1(_0584_),
    .A2(_0585_),
    .B(_0583_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1229_ (.A1(_0451_),
    .A2(_0580_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1230_ (.A1(\uart.divisor[14] ),
    .A2(_0575_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1231_ (.A1(_0586_),
    .A2(_0587_),
    .B(_0583_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1232_ (.A1(_0454_),
    .A2(_0580_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1233_ (.A1(\uart.divisor[15] ),
    .A2(_0575_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1234_ (.A1(_0588_),
    .A2(_0589_),
    .B(_0583_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1235_ (.A1(_0425_),
    .A2(_0476_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1236_ (.I(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1237_ (.I(_0590_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1238_ (.A1(\spi.divisor[0] ),
    .A2(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1239_ (.A1(_0280_),
    .A2(_0591_),
    .B(_0593_),
    .C(_0432_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1240_ (.A1(\spi.divisor[1] ),
    .A2(_0592_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1241_ (.A1(_0287_),
    .A2(_0591_),
    .B(_0594_),
    .C(_0432_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1242_ (.A1(_0425_),
    .A2(_0476_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1243_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1244_ (.A1(_0435_),
    .A2(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1245_ (.A1(_0256_),
    .A2(_0596_),
    .B(_0597_),
    .C(_0434_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1246_ (.A1(_0440_),
    .A2(_0596_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1247_ (.A1(_0251_),
    .A2(_0596_),
    .B(_0598_),
    .C(_0434_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1248_ (.A1(_0444_),
    .A2(_0595_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1249_ (.A1(\spi.divisor[4] ),
    .A2(_0591_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1250_ (.I(_0420_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1251_ (.A1(_0599_),
    .A2(_0600_),
    .B(_0601_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1252_ (.A1(_0448_),
    .A2(_0595_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1253_ (.A1(\spi.divisor[5] ),
    .A2(_0592_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1254_ (.A1(_0602_),
    .A2(_0603_),
    .B(_0601_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1255_ (.A1(_0451_),
    .A2(_0590_),
    .B(_0488_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1256_ (.A1(_0250_),
    .A2(_0591_),
    .B(_0604_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1257_ (.A1(_0454_),
    .A2(_0595_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1258_ (.A1(\spi.divisor[7] ),
    .A2(_0592_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1259_ (.A1(_0605_),
    .A2(_0606_),
    .B(_0601_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1260_ (.I(_0509_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1261_ (.I(\uart.receive_div_counter[0] ),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1262_ (.A1(\uart.receiving ),
    .A2(_0552_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1263_ (.I(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1264_ (.I(_0537_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1265_ (.I(_0548_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1266_ (.A1(_0611_),
    .A2(_0612_),
    .B(\uart.receiving ),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1267_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1268_ (.A1(_0608_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1269_ (.A1(_0608_),
    .A2(_0610_),
    .B(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1270_ (.A1(_0607_),
    .A2(_0616_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1271_ (.I(\uart.receive_div_counter[1] ),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1272_ (.A1(_0615_),
    .A2(_0610_),
    .B(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1273_ (.I(_0617_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1274_ (.A1(_0611_),
    .A2(_0612_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1275_ (.A1(_0551_),
    .A2(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1276_ (.I(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1277_ (.A1(_0619_),
    .A2(_0608_),
    .A3(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1278_ (.A1(_0618_),
    .A2(_0623_),
    .B(_0601_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1279_ (.I(\uart.receive_div_counter[2] ),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1280_ (.I(_0609_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1281_ (.A1(_0624_),
    .A2(_0617_),
    .A3(\uart.receive_div_counter[0] ),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1282_ (.I(_0621_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1283_ (.A1(_0624_),
    .A2(_0625_),
    .B1(_0626_),
    .B2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1284_ (.A1(_0617_),
    .A2(_0608_),
    .B(_0624_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1285_ (.A1(_0246_),
    .A2(_0628_),
    .A3(_0629_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1286_ (.I(\uart.receive_div_counter[3] ),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1287_ (.A1(\uart.receive_div_counter[3] ),
    .A2(_0625_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1288_ (.I(_0621_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1289_ (.A1(\uart.receive_div_counter[3] ),
    .A2(_0624_),
    .A3(\uart.receive_div_counter[1] ),
    .A4(\uart.receive_div_counter[0] ),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1290_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1291_ (.A1(_0632_),
    .A2(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1292_ (.I(_0245_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1293_ (.A1(_0630_),
    .A2(_0626_),
    .B1(_0631_),
    .B2(_0635_),
    .C(_0636_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1294_ (.I(\uart.receive_div_counter[4] ),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1295_ (.A1(_0637_),
    .A2(_0634_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1296_ (.A1(_0551_),
    .A2(net1),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1297_ (.A1(_0614_),
    .A2(_0638_),
    .B(_0639_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1298_ (.A1(\uart.receive_div_counter[4] ),
    .A2(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1299_ (.I(_0613_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1300_ (.A1(\uart.receive_div_counter[4] ),
    .A2(_0642_),
    .A3(_0634_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1301_ (.I(_0420_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1302_ (.A1(_0641_),
    .A2(_0643_),
    .B(_0644_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1303_ (.I(\uart.receive_div_counter[5] ),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1304_ (.A1(_0645_),
    .A2(_0637_),
    .A3(_0634_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1305_ (.A1(_0645_),
    .A2(_0640_),
    .B1(_0646_),
    .B2(_0622_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1306_ (.A1(_0607_),
    .A2(_0647_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1307_ (.A1(\uart.receive_div_counter[6] ),
    .A2(_0645_),
    .A3(_0638_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1308_ (.A1(_0614_),
    .A2(_0648_),
    .B(_0639_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1309_ (.A1(\uart.receive_div_counter[6] ),
    .A2(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1310_ (.A1(_0642_),
    .A2(_0648_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1311_ (.A1(_0645_),
    .A2(_0638_),
    .A3(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1312_ (.A1(_0650_),
    .A2(_0652_),
    .B(_0644_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1313_ (.A1(\uart.receive_div_counter[7] ),
    .A2(_0649_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1314_ (.I(\uart.receive_div_counter[7] ),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1315_ (.A1(_0654_),
    .A2(_0622_),
    .A3(_0648_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1316_ (.A1(_0653_),
    .A2(_0655_),
    .B(_0644_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1317_ (.A1(\uart.receive_div_counter[7] ),
    .A2(\uart.receive_div_counter[6] ),
    .A3(\uart.receive_div_counter[5] ),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1318_ (.A1(_0637_),
    .A2(_0633_),
    .A3(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1319_ (.I(\uart.receive_div_counter[8] ),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1320_ (.A1(_0658_),
    .A2(_0657_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1321_ (.A1(_0642_),
    .A2(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1322_ (.A1(_0614_),
    .A2(_0659_),
    .B(_0639_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1323_ (.A1(_0657_),
    .A2(_0660_),
    .B1(_0661_),
    .B2(_0658_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1324_ (.A1(_0607_),
    .A2(_0662_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1325_ (.I(\uart.receive_div_counter[9] ),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1326_ (.A1(_0663_),
    .A2(_0661_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1327_ (.I(_0663_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1328_ (.A1(_0665_),
    .A2(_0622_),
    .A3(_0659_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1329_ (.A1(_0664_),
    .A2(_0666_),
    .B(_0644_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1330_ (.A1(_0663_),
    .A2(_0658_),
    .A3(_0657_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1331_ (.A1(_0632_),
    .A2(_0667_),
    .B(\uart.receive_div_counter[10] ),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1332_ (.A1(\uart.receive_div_counter[10] ),
    .A2(_0667_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1333_ (.A1(_0627_),
    .A2(_0669_),
    .B(_0609_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1334_ (.A1(_0246_),
    .A2(_0668_),
    .A3(_0670_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1335_ (.I(\uart.receive_div_counter[11] ),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1336_ (.A1(_0642_),
    .A2(_0669_),
    .B(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1337_ (.A1(_0369_),
    .A2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1338_ (.A1(\uart.receive_div_counter[11] ),
    .A2(_0670_),
    .B(_0673_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1339_ (.A1(\uart.receive_div_counter[11] ),
    .A2(\uart.receive_div_counter[10] ),
    .A3(_0663_),
    .A4(_0658_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1340_ (.A1(_0637_),
    .A2(_0633_),
    .A3(_0656_),
    .A4(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1341_ (.I(\uart.receive_div_counter[12] ),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1342_ (.A1(_0676_),
    .A2(_0675_),
    .B(_0613_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1343_ (.A1(_0675_),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1344_ (.A1(_0625_),
    .A2(_0677_),
    .B(_0676_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1345_ (.I(_0419_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1346_ (.I(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1347_ (.A1(_0678_),
    .A2(_0679_),
    .B(_0681_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1348_ (.A1(_0625_),
    .A2(_0677_),
    .B(\uart.receive_div_counter[13] ),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1349_ (.I(\uart.receive_div_counter[13] ),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1350_ (.A1(_0683_),
    .A2(_0676_),
    .A3(_0632_),
    .A4(_0675_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1351_ (.A1(_0682_),
    .A2(_0684_),
    .B(_0681_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1352_ (.I(\uart.receive_div_counter[14] ),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1353_ (.A1(\uart.receive_div_counter[13] ),
    .A2(_0676_),
    .A3(_0675_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1354_ (.A1(_0685_),
    .A2(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1355_ (.A1(_0685_),
    .A2(_0686_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1356_ (.A1(_0632_),
    .A2(_0687_),
    .A3(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1357_ (.A1(_0685_),
    .A2(_0610_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1358_ (.A1(_0689_),
    .A2(_0690_),
    .B(_0681_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1359_ (.I(\uart.receive_div_counter[15] ),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1360_ (.A1(_0685_),
    .A2(_0627_),
    .A3(_0686_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1361_ (.A1(_0627_),
    .A2(_0688_),
    .B(_0609_),
    .C(_0691_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1362_ (.I(_0353_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1363_ (.A1(_0691_),
    .A2(_0692_),
    .B(_0693_),
    .C(_0694_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1364_ (.A1(\uart.receive_counter[3] ),
    .A2(_0562_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1365_ (.A1(_0611_),
    .A2(_0612_),
    .A3(_0695_),
    .B(\uart.receiving ),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1366_ (.A1(_0639_),
    .A2(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1367_ (.I(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1368_ (.A1(_0551_),
    .A2(_0611_),
    .A3(_0612_),
    .A4(_0695_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1369_ (.I(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1370_ (.A1(\uart.receive_buff[0] ),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\uart.receive_buff[1] ),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1371_ (.A1(_0607_),
    .A2(_0701_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1372_ (.I(_0509_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1373_ (.A1(\uart.receive_buff[1] ),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\uart.receive_buff[2] ),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1374_ (.A1(_0702_),
    .A2(_0703_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1375_ (.A1(\uart.receive_buff[2] ),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\uart.receive_buff[3] ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1376_ (.A1(_0702_),
    .A2(_0704_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1377_ (.I(_0699_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1378_ (.A1(\uart.receive_buff[3] ),
    .A2(_0698_),
    .B1(_0705_),
    .B2(\uart.receive_buff[4] ),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1379_ (.A1(_0702_),
    .A2(_0706_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1380_ (.A1(\uart.receive_buff[4] ),
    .A2(_0697_),
    .B1(_0705_),
    .B2(\uart.receive_buff[5] ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1381_ (.A1(_0702_),
    .A2(_0707_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1382_ (.I(_0509_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1383_ (.A1(\uart.receive_buff[5] ),
    .A2(_0697_),
    .B1(_0705_),
    .B2(\uart.receive_buff[6] ),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1384_ (.A1(_0708_),
    .A2(_0709_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1385_ (.A1(\uart.receive_buff[6] ),
    .A2(_0697_),
    .B1(_0705_),
    .B2(\uart.receive_buff[7] ),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1386_ (.A1(_0708_),
    .A2(_0710_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1387_ (.A1(\uart.receive_buff[7] ),
    .A2(_0700_),
    .B(_0431_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1388_ (.A1(_0552_),
    .A2(_0696_),
    .B(_0711_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1389_ (.A1(_0526_),
    .A2(_0537_),
    .A3(_0548_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1390_ (.A1(_0712_),
    .A2(_0695_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1391_ (.I(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1392_ (.A1(_0246_),
    .A2(_0610_),
    .A3(_0714_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1393_ (.I(\uart.div_counter[15] ),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1394_ (.A1(_0715_),
    .A2(\uart.divisor[15] ),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1395_ (.A1(\uart.div_counter[2] ),
    .A2(\uart.divisor[2] ),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1396_ (.A1(\uart.div_counter[11] ),
    .A2(\uart.divisor[11] ),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1397_ (.A1(\uart.div_counter[6] ),
    .A2(\uart.divisor[6] ),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1398_ (.A1(_0718_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1399_ (.A1(\uart.div_counter[13] ),
    .A2(\uart.divisor[13] ),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1400_ (.A1(\uart.div_counter[4] ),
    .A2(\uart.divisor[4] ),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1401_ (.A1(\uart.div_counter[5] ),
    .A2(\uart.divisor[5] ),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1402_ (.A1(\uart.div_counter[7] ),
    .A2(\uart.divisor[7] ),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1403_ (.A1(_0721_),
    .A2(_0722_),
    .A3(_0723_),
    .A4(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _1404_ (.A1(_0716_),
    .A2(_0717_),
    .A3(_0720_),
    .A4(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1405_ (.I(_0726_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1406_ (.A1(\uart.div_counter[9] ),
    .A2(\uart.divisor[9] ),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1407_ (.A1(\uart.div_counter[1] ),
    .A2(\uart.divisor[1] ),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1408_ (.A1(\uart.div_counter[3] ),
    .A2(\uart.divisor[3] ),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1409_ (.A1(\uart.div_counter[12] ),
    .A2(\uart.divisor[12] ),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1410_ (.A1(_0728_),
    .A2(_0729_),
    .A3(_0730_),
    .A4(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1411_ (.A1(\uart.div_counter[14] ),
    .A2(\uart.divisor[14] ),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1412_ (.A1(\uart.div_counter[10] ),
    .A2(\uart.divisor[10] ),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1413_ (.A1(\uart.div_counter[8] ),
    .A2(\uart.divisor[8] ),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1414_ (.A1(\uart.div_counter[0] ),
    .A2(\uart.divisor[0] ),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1415_ (.A1(_0733_),
    .A2(_0734_),
    .A3(_0735_),
    .A4(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1416_ (.A1(_0732_),
    .A2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1417_ (.I(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1418_ (.I(\uart.counter[0] ),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1419_ (.A1(\uart.busy ),
    .A2(_0275_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1420_ (.A1(_0474_),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1421_ (.A1(_0740_),
    .A2(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1422_ (.A1(_0727_),
    .A2(_0739_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1423_ (.A1(\uart.counter[0] ),
    .A2(\uart.counter[1] ),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1424_ (.A1(\uart.counter[3] ),
    .A2(\uart.counter[2] ),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1425_ (.A1(_0745_),
    .A2(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1426_ (.I(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1427_ (.A1(_0419_),
    .A2(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1428_ (.I(_0749_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1429_ (.A1(_0726_),
    .A2(_0738_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1430_ (.A1(_0740_),
    .A2(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1431_ (.A1(_0744_),
    .A2(_0126_),
    .A3(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1432_ (.I(_0752_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1433_ (.I(\uart.counter[1] ),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1434_ (.A1(_0475_),
    .A2(_0741_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1435_ (.I(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1436_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1437_ (.A1(_0727_),
    .A2(_0739_),
    .A3(_0746_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1438_ (.A1(_0756_),
    .A2(_0757_),
    .B(_0751_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1439_ (.A1(_0740_),
    .A2(_0753_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1440_ (.I(_0750_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1441_ (.A1(_0753_),
    .A2(_0758_),
    .B1(_0759_),
    .B2(_0760_),
    .C(_0636_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1442_ (.A1(\uart.counter[2] ),
    .A2(_0745_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1443_ (.A1(_0760_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1444_ (.I(_0742_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1445_ (.A1(_0727_),
    .A2(_0739_),
    .B(_0763_),
    .C(\uart.counter[2] ),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1446_ (.A1(_0762_),
    .A2(_0764_),
    .B(_0636_),
    .C(_0748_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1447_ (.I(\uart.counter[3] ),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1448_ (.A1(_0740_),
    .A2(\uart.counter[1] ),
    .A3(\uart.counter[2] ),
    .B(\uart.counter[3] ),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1449_ (.A1(_0726_),
    .A2(_0738_),
    .A3(_0747_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1450_ (.I(_0767_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1451_ (.I(_0768_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1452_ (.A1(_0765_),
    .A2(_0763_),
    .B1(_0766_),
    .B2(_0769_),
    .C(_0357_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1453_ (.A1(\uart.data_buff[1] ),
    .A2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1454_ (.I(\uart.data_buff[0] ),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1455_ (.I(_0768_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1456_ (.A1(_0771_),
    .A2(_0756_),
    .A3(_0772_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1457_ (.A1(_0770_),
    .A2(_0773_),
    .B(_0681_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1458_ (.I(\uart.data_buff[2] ),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1459_ (.I(_0769_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1460_ (.A1(_0279_),
    .A2(_0742_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1461_ (.A1(\uart.data_buff[1] ),
    .A2(_0763_),
    .B(_0772_),
    .C(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1462_ (.A1(_0774_),
    .A2(_0775_),
    .B(_0777_),
    .C(_0694_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1463_ (.I(\uart.data_buff[3] ),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1464_ (.I(_0754_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1465_ (.A1(_0774_),
    .A2(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1466_ (.A1(net8),
    .A2(_0756_),
    .B(_0772_),
    .C(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1467_ (.A1(_0778_),
    .A2(_0775_),
    .B(_0781_),
    .C(_0694_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1468_ (.I(\uart.data_buff[4] ),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1469_ (.I(_0767_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1470_ (.A1(_0778_),
    .A2(_0779_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1471_ (.A1(_0435_),
    .A2(_0756_),
    .B(_0783_),
    .C(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1472_ (.A1(_0782_),
    .A2(_0775_),
    .B(_0785_),
    .C(_0694_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1473_ (.I(\uart.data_buff[5] ),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1474_ (.I(_0755_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1475_ (.A1(_0782_),
    .A2(_0779_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1476_ (.A1(_0440_),
    .A2(_0787_),
    .B(_0783_),
    .C(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1477_ (.I(_0245_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1478_ (.A1(_0786_),
    .A2(_0775_),
    .B(_0789_),
    .C(_0790_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1479_ (.I(\uart.data_buff[6] ),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1480_ (.I(_0772_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1481_ (.I(_0755_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1482_ (.A1(_0786_),
    .A2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1483_ (.A1(_0444_),
    .A2(_0787_),
    .B(_0783_),
    .C(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1484_ (.A1(_0791_),
    .A2(_0792_),
    .B(_0795_),
    .C(_0790_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1485_ (.I(\uart.data_buff[7] ),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1486_ (.A1(_0791_),
    .A2(_0793_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1487_ (.A1(_0448_),
    .A2(_0787_),
    .B(_0783_),
    .C(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1488_ (.A1(_0796_),
    .A2(_0792_),
    .B(_0798_),
    .C(_0790_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1489_ (.I(\uart.data_buff[8] ),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1490_ (.A1(_0796_),
    .A2(_0793_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1491_ (.A1(_0451_),
    .A2(_0787_),
    .B(_0768_),
    .C(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1492_ (.A1(_0799_),
    .A2(_0792_),
    .B(_0801_),
    .C(_0790_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1493_ (.I(\uart.data_buff[9] ),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1494_ (.A1(_0799_),
    .A2(_0793_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1495_ (.A1(_0454_),
    .A2(_0779_),
    .B(_0768_),
    .C(_0803_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1496_ (.I(_0245_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1497_ (.A1(_0802_),
    .A2(_0792_),
    .B(_0804_),
    .C(_0805_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1498_ (.A1(_0802_),
    .A2(_0763_),
    .B(_0769_),
    .C(_0805_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1499_ (.I(\uart.div_counter[0] ),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1500_ (.A1(_0745_),
    .A2(_0746_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1501_ (.A1(_0755_),
    .A2(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1502_ (.I(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1503_ (.A1(_0727_),
    .A2(_0739_),
    .B(_0807_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1504_ (.I(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1505_ (.A1(_0806_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1506_ (.A1(_0806_),
    .A2(_0809_),
    .B(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1507_ (.A1(_0708_),
    .A2(_0813_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1508_ (.I(\uart.div_counter[1] ),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1509_ (.A1(_0812_),
    .A2(_0809_),
    .B(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1510_ (.I(_0814_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1511_ (.A1(_0750_),
    .A2(_0748_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1512_ (.I(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1513_ (.A1(_0816_),
    .A2(_0806_),
    .A3(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1514_ (.I(_0680_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1515_ (.A1(_0815_),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1516_ (.I(\uart.div_counter[2] ),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1517_ (.A1(_0821_),
    .A2(_0814_),
    .A3(\uart.div_counter[0] ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1518_ (.I(_0817_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1519_ (.A1(_0821_),
    .A2(_0809_),
    .B1(_0822_),
    .B2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1520_ (.A1(_0814_),
    .A2(_0806_),
    .B(_0821_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1521_ (.A1(_0636_),
    .A2(_0824_),
    .A3(_0825_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1522_ (.I(\uart.div_counter[3] ),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1523_ (.A1(\uart.div_counter[3] ),
    .A2(_0821_),
    .A3(\uart.div_counter[1] ),
    .A4(\uart.div_counter[0] ),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1524_ (.I(_0144_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1525_ (.A1(\uart.div_counter[3] ),
    .A2(_0808_),
    .B1(_0145_),
    .B2(_0823_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1526_ (.A1(_0826_),
    .A2(_0822_),
    .B(_0146_),
    .C(_0805_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1527_ (.I(\uart.div_counter[4] ),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1528_ (.A1(_0147_),
    .A2(_0145_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1529_ (.A1(_0742_),
    .A2(_0748_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1530_ (.A1(_0811_),
    .A2(_0148_),
    .B(_0149_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1531_ (.A1(\uart.div_counter[4] ),
    .A2(_0150_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1532_ (.I(_0810_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1533_ (.A1(\uart.div_counter[4] ),
    .A2(_0152_),
    .A3(_0145_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1534_ (.A1(_0151_),
    .A2(_0153_),
    .B(_0820_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1535_ (.I(\uart.div_counter[5] ),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1536_ (.A1(_0154_),
    .A2(_0147_),
    .A3(_0145_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1537_ (.A1(_0154_),
    .A2(_0150_),
    .B1(_0155_),
    .B2(_0818_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1538_ (.A1(_0708_),
    .A2(_0156_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1539_ (.I(_0810_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1540_ (.A1(\uart.div_counter[6] ),
    .A2(_0154_),
    .A3(_0148_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1541_ (.I(_0149_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1542_ (.A1(_0157_),
    .A2(_0158_),
    .B(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1543_ (.A1(\uart.div_counter[6] ),
    .A2(_0160_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1544_ (.A1(_0152_),
    .A2(_0158_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1545_ (.A1(_0154_),
    .A2(_0148_),
    .A3(_0162_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1546_ (.A1(_0161_),
    .A2(_0163_),
    .B(_0820_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1547_ (.A1(\uart.div_counter[7] ),
    .A2(_0160_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1548_ (.I(\uart.div_counter[7] ),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1549_ (.A1(_0165_),
    .A2(_0818_),
    .A3(_0158_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1550_ (.A1(_0164_),
    .A2(_0166_),
    .B(_0820_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1551_ (.I(_0390_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1552_ (.A1(\uart.div_counter[7] ),
    .A2(\uart.div_counter[6] ),
    .A3(\uart.div_counter[5] ),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1553_ (.A1(_0147_),
    .A2(_0144_),
    .A3(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1554_ (.A1(\uart.div_counter[8] ),
    .A2(_0169_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1555_ (.I(_0170_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1556_ (.A1(_0157_),
    .A2(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1557_ (.A1(_0811_),
    .A2(_0171_),
    .B(_0159_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1558_ (.A1(_0169_),
    .A2(_0172_),
    .B1(_0173_),
    .B2(\uart.div_counter[8] ),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1559_ (.A1(_0167_),
    .A2(_0174_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1560_ (.I(\uart.div_counter[9] ),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1561_ (.A1(_0175_),
    .A2(_0173_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1562_ (.I(_0175_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1563_ (.A1(_0177_),
    .A2(_0818_),
    .A3(_0171_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1564_ (.I(_0680_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1565_ (.A1(_0176_),
    .A2(_0178_),
    .B(_0179_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1566_ (.A1(\uart.div_counter[10] ),
    .A2(_0175_),
    .A3(_0170_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1567_ (.A1(_0811_),
    .A2(_0180_),
    .B(_0159_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1568_ (.A1(\uart.div_counter[10] ),
    .A2(_0181_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1569_ (.A1(_0157_),
    .A2(_0180_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1570_ (.A1(_0175_),
    .A2(_0171_),
    .A3(_0183_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1571_ (.A1(_0182_),
    .A2(_0184_),
    .B(_0179_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1572_ (.A1(\uart.div_counter[11] ),
    .A2(_0152_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1573_ (.A1(_0180_),
    .A2(_0185_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1574_ (.A1(\uart.div_counter[11] ),
    .A2(_0181_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1575_ (.A1(_0186_),
    .A2(_0187_),
    .B(_0179_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1576_ (.I(\uart.div_counter[12] ),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1577_ (.I(_0188_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1578_ (.A1(\uart.div_counter[11] ),
    .A2(\uart.div_counter[10] ),
    .A3(\uart.div_counter[9] ),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1579_ (.A1(\uart.div_counter[8] ),
    .A2(_0169_),
    .A3(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1580_ (.A1(_0189_),
    .A2(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1581_ (.A1(_0810_),
    .A2(_0192_),
    .B(_0149_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1582_ (.A1(_0188_),
    .A2(_0157_),
    .A3(_0191_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1583_ (.A1(_0188_),
    .A2(_0193_),
    .B(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1584_ (.A1(_0167_),
    .A2(_0195_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1585_ (.A1(\uart.div_counter[13] ),
    .A2(_0152_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1586_ (.A1(\uart.div_counter[13] ),
    .A2(_0193_),
    .B1(_0196_),
    .B2(_0192_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1587_ (.A1(_0167_),
    .A2(_0197_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1588_ (.I(\uart.div_counter[14] ),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1589_ (.A1(\uart.div_counter[13] ),
    .A2(_0188_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1590_ (.A1(_0198_),
    .A2(_0191_),
    .A3(_0199_),
    .B(_0817_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1591_ (.A1(_0191_),
    .A2(_0199_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1592_ (.A1(_0823_),
    .A2(_0201_),
    .B(\uart.div_counter[14] ),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1593_ (.A1(_0159_),
    .A2(_0200_),
    .B(_0202_),
    .C(_0805_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1594_ (.A1(_0715_),
    .A2(_0809_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1595_ (.A1(\uart.div_counter[14] ),
    .A2(_0823_),
    .A3(_0201_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1596_ (.A1(_0200_),
    .A2(_0203_),
    .B1(_0204_),
    .B2(_0715_),
    .C(_0357_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1597_ (.A1(_0712_),
    .A2(_0695_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1598_ (.I(_0205_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1599_ (.A1(net8),
    .A2(_0566_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1600_ (.A1(\uart.has_byte ),
    .A2(_0207_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1601_ (.A1(_0206_),
    .A2(_0208_),
    .B(_0179_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1602_ (.I(net15),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1603_ (.A1(_0276_),
    .A2(_0394_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1604_ (.I(_0210_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1605_ (.A1(_0209_),
    .A2(_0396_),
    .B1(_0211_),
    .B2(_0399_),
    .C(_0357_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1606_ (.A1(\spi.data_in_buff[0] ),
    .A2(_0396_),
    .B1(_0211_),
    .B2(\spi.data_in_buff[1] ),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1607_ (.A1(_0167_),
    .A2(_0212_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1608_ (.I(_0390_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1609_ (.I(_0395_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1610_ (.A1(\spi.data_in_buff[1] ),
    .A2(_0214_),
    .B1(_0211_),
    .B2(\spi.data_in_buff[2] ),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1611_ (.A1(_0213_),
    .A2(_0215_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1612_ (.A1(\spi.data_in_buff[2] ),
    .A2(_0214_),
    .B1(_0211_),
    .B2(\spi.data_in_buff[3] ),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1613_ (.A1(_0213_),
    .A2(_0216_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1614_ (.I(_0210_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1615_ (.A1(\spi.data_in_buff[3] ),
    .A2(_0214_),
    .B1(_0217_),
    .B2(\spi.data_in_buff[4] ),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1616_ (.A1(_0213_),
    .A2(_0218_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1617_ (.A1(\spi.data_in_buff[4] ),
    .A2(_0214_),
    .B1(_0217_),
    .B2(\spi.data_in_buff[5] ),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1618_ (.A1(_0213_),
    .A2(_0219_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1619_ (.A1(\spi.data_in_buff[5] ),
    .A2(_0395_),
    .B1(_0217_),
    .B2(\spi.data_in_buff[6] ),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1620_ (.A1(_0354_),
    .A2(_0220_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1621_ (.A1(\spi.data_in_buff[6] ),
    .A2(_0395_),
    .B1(_0217_),
    .B2(\spi.data_in_buff[7] ),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1622_ (.A1(_0354_),
    .A2(_0221_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1623_ (.A1(_0771_),
    .A2(_0760_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1624_ (.A1(net17),
    .A2(_0760_),
    .B(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1625_ (.A1(_0126_),
    .A2(_0223_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1626_ (.A1(\uart.receive_buff[0] ),
    .A2(_0714_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1627_ (.A1(\uart.dout[0] ),
    .A2(_0206_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1628_ (.I(_0680_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1629_ (.A1(_0224_),
    .A2(_0225_),
    .B(_0226_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1630_ (.A1(\uart.receive_buff[1] ),
    .A2(_0714_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1631_ (.A1(\uart.dout[1] ),
    .A2(_0206_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1632_ (.A1(_0227_),
    .A2(_0228_),
    .B(_0226_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1633_ (.A1(\uart.receive_buff[2] ),
    .A2(_0714_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1634_ (.A1(\uart.dout[2] ),
    .A2(_0206_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1635_ (.A1(_0229_),
    .A2(_0230_),
    .B(_0226_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1636_ (.I(_0713_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1637_ (.A1(\uart.receive_buff[3] ),
    .A2(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1638_ (.I(_0205_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1639_ (.A1(\uart.dout[3] ),
    .A2(_0233_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1640_ (.A1(_0232_),
    .A2(_0234_),
    .B(_0226_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1641_ (.A1(\uart.receive_buff[4] ),
    .A2(_0231_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1642_ (.A1(\uart.dout[4] ),
    .A2(_0233_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1643_ (.I(_0353_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1644_ (.A1(_0235_),
    .A2(_0236_),
    .B(_0237_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1645_ (.A1(\uart.receive_buff[5] ),
    .A2(_0231_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1646_ (.A1(\uart.dout[5] ),
    .A2(_0233_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1647_ (.A1(_0238_),
    .A2(_0239_),
    .B(_0237_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1648_ (.A1(\uart.receive_buff[6] ),
    .A2(_0231_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1649_ (.A1(\uart.dout[6] ),
    .A2(_0233_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1650_ (.A1(_0240_),
    .A2(_0241_),
    .B(_0237_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1651_ (.A1(\uart.receive_buff[7] ),
    .A2(_0713_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1652_ (.A1(\uart.dout[7] ),
    .A2(_0205_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1653_ (.A1(_0242_),
    .A2(_0243_),
    .B(_0237_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1654_ (.D(_0000_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(\spi.data_out_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1655_ (.D(_0001_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.data_out_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1656_ (.D(_0002_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.data_out_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1657_ (.D(_0003_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.data_out_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1658_ (.D(_0004_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.data_out_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1659_ (.D(_0005_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(\spi.data_out_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1660_ (.D(_0006_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(\spi.data_out_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1661_ (.D(_0007_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(\spi.data_out_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1662_ (.D(_0008_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1663_ (.D(_0009_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1664_ (.D(_0010_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1665_ (.D(_0011_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(\spi.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1666_ (.D(_0012_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\spi.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1667_ (.D(_0013_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.busy ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1668_ (.D(_0014_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.div_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1669_ (.D(_0015_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.div_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1670_ (.D(_0016_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.div_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1671_ (.D(_0017_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(\spi.div_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1672_ (.D(_0018_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(\spi.div_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1673_ (.D(_0019_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(\spi.div_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1674_ (.D(_0020_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(\spi.div_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1675_ (.D(_0021_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(\spi.div_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1676_ (.D(_0022_),
    .CLK(clknet_4_8_0_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1677_ (.D(_0023_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.dout[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1678_ (.D(_0024_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1679_ (.D(_0025_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.dout[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1680_ (.D(_0026_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.dout[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1681_ (.D(_0027_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.dout[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1682_ (.D(_0028_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1683_ (.D(_0029_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1684_ (.D(_0030_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1685_ (.D(_0031_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1686_ (.D(_0032_),
    .CLK(clknet_4_9_0_wb_clk_i),
    .Q(\uart.divisor[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1687_ (.D(_0033_),
    .CLK(clknet_4_9_0_wb_clk_i),
    .Q(\uart.divisor[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1688_ (.D(_0034_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.divisor[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1689_ (.D(_0035_),
    .CLK(clknet_4_9_0_wb_clk_i),
    .Q(\uart.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1690_ (.D(_0036_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1691_ (.D(_0037_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.divisor[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1692_ (.D(_0038_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1693_ (.D(_0039_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1694_ (.D(_0040_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1695_ (.D(_0041_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1696_ (.D(_0042_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1697_ (.D(_0043_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1698_ (.D(_0044_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1699_ (.D(_0045_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1700_ (.D(_0046_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1701_ (.D(_0047_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1702_ (.D(_0048_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1703_ (.D(_0049_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\uart.receive_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1704_ (.D(_0050_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\uart.receive_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1705_ (.D(_0051_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\uart.receive_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1706_ (.D(_0052_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\uart.receive_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1707_ (.D(_0053_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(uart_ien));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1708_ (.D(_0054_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\uart.divisor[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1709_ (.D(_0055_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\uart.divisor[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1710_ (.D(_0056_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.divisor[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1711_ (.D(_0057_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.divisor[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1712_ (.D(_0058_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\uart.divisor[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1713_ (.D(_0059_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.divisor[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1714_ (.D(_0060_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\uart.divisor[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1715_ (.D(_0061_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\uart.divisor[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1716_ (.D(_0062_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.divisor[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1717_ (.D(_0063_),
    .CLK(clknet_4_9_0_wb_clk_i),
    .Q(\spi.divisor[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1718_ (.D(_0064_),
    .CLK(clknet_4_9_0_wb_clk_i),
    .Q(\spi.divisor[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1719_ (.D(_0065_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\spi.divisor[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1720_ (.D(_0066_),
    .CLK(clknet_4_9_0_wb_clk_i),
    .Q(\spi.divisor[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1721_ (.D(_0067_),
    .CLK(clknet_4_9_0_wb_clk_i),
    .Q(\spi.divisor[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1722_ (.D(_0068_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(\spi.divisor[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1723_ (.D(_0069_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(\spi.divisor[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1724_ (.D(_0070_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.receive_div_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1725_ (.D(_0071_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1726_ (.D(_0072_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1727_ (.D(_0073_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1728_ (.D(_0074_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1729_ (.D(_0075_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receive_div_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1730_ (.D(_0076_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receive_div_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1731_ (.D(_0077_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receive_div_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1732_ (.D(_0078_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receive_div_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1733_ (.D(_0079_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1734_ (.D(_0080_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1735_ (.D(_0081_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1736_ (.D(_0082_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\uart.receive_div_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1737_ (.D(_0083_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\uart.receive_div_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1738_ (.D(_0084_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\uart.receive_div_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1739_ (.D(_0085_),
    .CLK(clknet_4_7_0_wb_clk_i),
    .Q(\uart.receive_div_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1740_ (.D(_0086_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receive_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1741_ (.D(_0087_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receive_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1742_ (.D(_0088_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\uart.receive_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1743_ (.D(_0089_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\uart.receive_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1744_ (.D(_0090_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\uart.receive_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1745_ (.D(_0091_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\uart.receive_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1746_ (.D(_0092_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\uart.receive_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1747_ (.D(_0093_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receive_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1748_ (.D(_0094_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\uart.receiving ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1749_ (.D(_0095_),
    .CLK(clknet_4_1_0_wb_clk_i),
    .Q(\uart.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1750_ (.D(_0096_),
    .CLK(clknet_4_1_0_wb_clk_i),
    .Q(\uart.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1751_ (.D(_0097_),
    .CLK(clknet_4_1_0_wb_clk_i),
    .Q(\uart.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1752_ (.D(_0098_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\uart.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1753_ (.D(_0099_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\uart.data_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1754_ (.D(_0100_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\uart.data_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1755_ (.D(_0101_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\uart.data_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1756_ (.D(_0102_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\uart.data_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1757_ (.D(_0103_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\uart.data_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1758_ (.D(_0104_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\uart.data_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1759_ (.D(_0105_),
    .CLK(clknet_4_3_0_wb_clk_i),
    .Q(\uart.data_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1760_ (.D(_0106_),
    .CLK(clknet_4_1_0_wb_clk_i),
    .Q(\uart.data_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1761_ (.D(_0107_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\uart.data_buff[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1762_ (.D(_0108_),
    .CLK(clknet_4_1_0_wb_clk_i),
    .Q(\uart.data_buff[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1763_ (.D(_0109_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\uart.div_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1764_ (.D(_0110_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1765_ (.D(_0111_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\uart.div_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1766_ (.D(_0112_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\uart.div_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1767_ (.D(_0113_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\uart.div_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1768_ (.D(_0114_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\uart.div_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1769_ (.D(_0115_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\uart.div_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1770_ (.D(_0116_),
    .CLK(clknet_4_5_0_wb_clk_i),
    .Q(\uart.div_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1771_ (.D(_0117_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1772_ (.D(_0118_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1773_ (.D(_0119_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1774_ (.D(_0120_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1775_ (.D(_0121_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1776_ (.D(_0122_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1777_ (.D(_0123_),
    .CLK(clknet_4_4_0_wb_clk_i),
    .Q(\uart.div_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1778_ (.D(_0124_),
    .CLK(clknet_4_6_0_wb_clk_i),
    .Q(\uart.div_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1779_ (.D(_0125_),
    .CLK(clknet_4_11_0_wb_clk_i),
    .Q(\uart.has_byte ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1780_ (.D(_0126_),
    .CLK(clknet_4_1_0_wb_clk_i),
    .Q(\uart.busy ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1781_ (.D(_0127_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.data_in_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1782_ (.D(_0128_),
    .CLK(clknet_4_1_0_wb_clk_i),
    .Q(\spi.data_in_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1783_ (.D(_0129_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\spi.data_in_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1784_ (.D(_0130_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\spi.data_in_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1785_ (.D(_0131_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\spi.data_in_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1786_ (.D(_0132_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\spi.data_in_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1787_ (.D(_0133_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.data_in_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1788_ (.D(_0134_),
    .CLK(clknet_4_2_0_wb_clk_i),
    .Q(\spi.data_in_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1789_ (.D(_0135_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1790_ (.D(_0136_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.dout[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1791_ (.D(_0137_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.dout[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1792_ (.D(_0138_),
    .CLK(clknet_4_12_0_wb_clk_i),
    .Q(\uart.dout[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1793_ (.D(_0139_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\uart.dout[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1794_ (.D(_0140_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\uart.dout[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1795_ (.D(_0141_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\uart.dout[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1796_ (.D(_0142_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\uart.dout[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1797_ (.D(_0143_),
    .CLK(clknet_4_14_0_wb_clk_i),
    .Q(\uart.dout[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1 (.I(RXD),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(data_in[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(data_in[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(data_in[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(data_in[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(data_in[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(io_in),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(rst),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(addr[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input3 (.I(addr[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(addr[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(bus_cyc),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(bus_we),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(data_in[0]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input8 (.I(data_in[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(data_in[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(TXD));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(irq3));
 gf180mcu_fd_sc_mcu7t5v0__tiel serial_ports_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel serial_ports_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel serial_ports_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tieh serial_ports_32 (.Z(net32));
 assign io_oeb[0] = net29;
 assign io_oeb[1] = net30;
 assign io_oeb[2] = net32;
 assign io_out[2] = net31;
endmodule

