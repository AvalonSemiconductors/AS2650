* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i wb_rst_i
XFILLER_79_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6209__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3691__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5968__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6914_ _1729_ _1818_ _2892_ _2895_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6845_ _0964_ _1109_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6776_ _2498_ _2757_ _2762_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3988_ _3297_ _3204_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6932__A3 _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5727_ _1040_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3746__A3 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6145__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5658_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4609_ _0626_ _0793_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _3251_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7328_ _0151_ clknet_3_3_0_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6448__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7259_ _0082_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3959__I _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6384__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6136__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6136__B2 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__A2 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5498__I0 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4960_ _0338_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3911_ _3258_ _3282_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4891_ _1009_ _1021_ _1031_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _2597_ _2612_ _2620_ _1600_ _1154_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3842_ _3353_ _3362_ _3377_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5178__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6561_ _2494_ _0583_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3773_ _3297_ _3299_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5512_ _1108_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6127__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _1098_ _1118_ _2501_ _1121_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5443_ _1045_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5374_ _1440_ _1441_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_99_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7113_ as2650.overflow _3065_ _0884_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _0499_ _3005_ _3008_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4256_ _0458_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4187_ _3393_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3664__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6828_ _1126_ _2684_ _2811_ _2812_ _2458_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6759_ _2613_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7427__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7094__A2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6774__B _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__C _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5580__A2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__C as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__I _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4110_ as2650.addr_buff\[7\] _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7085__A2 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5090_ as2650.stack\[5\]\[11\] _1247_ _1238_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4041_ _3324_ _3362_ _3574_ _3380_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5635__A3 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4843__A1 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6140__S0 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5992_ _0711_ _0921_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4943_ _0807_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4874_ _3208_ _3259_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _1419_ _2601_ _2603_ _1597_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3825_ _3360_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6544_ _2544_ _2545_ _2546_ _2550_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3756_ as2650.r123\[0\]\[0\] as2650.r123\[2\]\[0\] as2650.r123_2\[0\]\[0\] as2650.r123_2\[2\]\[0\]
+ _3125_ _3288_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_101_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5571__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6475_ _1652_ _2462_ _2484_ _2485_ _1095_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3687_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5426_ _1485_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4126__A3 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6520__A1 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5357_ _0925_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4308_ _0508_ _0510_ _3579_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7076__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5288_ as2650.stack\[0\]\[11\] _1377_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4893__I as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _3285_ _0798_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6823__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4239_ _3426_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6339__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5011__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3972__I _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7067__A2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4825__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4053__A2 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3610_ _3145_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4590_ _0772_ _0727_ _0776_ _0635_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4978__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__C _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1134_ _3341_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6502__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _0945_ _1328_ _1332_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6191_ as2650.pc\[6\] _1229_ _2130_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _0951_ _1276_ _1281_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7058__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6805__A2 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5073_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3619__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4024_ as2650.r0\[3\] _3331_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6861__C _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__B2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7272__CLK clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _0711_ _1739_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4044__A2 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4926_ _3165_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5792__A2 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _3146_ _3402_ _3256_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _3343_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5544__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6741__A1 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4888__I _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6527_ _1541_ _2522_ _1634_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3792__I _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3739_ _3274_ _3248_ _3189_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_109_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6458_ as2650.psu\[0\] _2469_ _1114_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5409_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6389_ _1300_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5512__I _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5480__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4283__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5668__B _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3967__I _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3794__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5535__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4798__I as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__A1 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__C _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7295__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6962__B _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4038__I _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5578__B _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5074__I1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5760_ _1423_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5774__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4711_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5691_ _0536_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7430_ _0253_ clknet_leaf_17_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4642_ _3252_ _3271_ _3466_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_129_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _0184_ clknet_leaf_54_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4573_ _0488_ _0760_ _0712_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _2250_ _2326_ _2327_ _2299_ _1981_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7292_ _0115_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6243_ _2258_ _2256_ _2257_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_104_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6856__C _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _1322_ _2059_ _2060_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ as2650.stack\[4\]\[11\] _1247_ _1266_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ _0947_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5462__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4265__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ _3437_ _3360_ _3502_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__5462__B2 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A2 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3787__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6962__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ _1888_ _1938_ _1980_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5765__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3776__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4909_ _3259_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5889_ _1487_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6714__B2 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4008__A2 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5756__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6801__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4192__A1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4247__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4991__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6930_ _2905_ _2906_ _2907_ _2910_ _1535_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _2687_ _2843_ _2844_ _1826_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ as2650.cycle\[5\] _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6792_ _0760_ _0467_ _2777_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5747__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3758__A1 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5743_ _1737_ _0621_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7310__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5674_ _1534_ _0822_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7413_ _0236_ clknet_leaf_24_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _0640_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4183__A1 _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _0167_ clknet_leaf_11_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4556_ _0741_ _0691_ _0744_ _0635_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3930__A1 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ _0098_ clknet_leaf_67_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4487_ _0675_ _0679_ _0649_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__7121__A1 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6226_ _2159_ _2238_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__A2 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5062__I _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _1260_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6088_ _1782_ _2100_ _2108_ _2008_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5039_ _0888_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5986__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5738__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__B2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6621__I _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5237__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4174__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5910__A2 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3921__A1 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5681__B _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput20 net20 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__A1 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput31 net31 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6496__C _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__S1 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5674__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5700__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__B _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7333__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__B _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4401__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6154__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4410_ as2650.r123\[1\]\[0\] _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4165__A1 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5390_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5901__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _3345_ _3572_ _0543_ _3323_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4986__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3890__I _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7103__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7060_ _1060_ _3019_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _3138_ as2650.r123\[0\]\[6\] _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6011_ _1440_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5417__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5968__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3979__A1 _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _2302_ _2893_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6844_ net35 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6917__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6775_ _1226_ _2700_ _2761_ _2699_ _1755_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3987_ _3383_ _3492_ _3520_ _3521_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _1499_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5657_ _0409_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4156__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _0583_ _0703_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4156__B2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5588_ _0875_ _1634_ _1018_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7327_ _0150_ clknet_leaf_3_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4539_ _0334_ _0712_ _0692_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _0081_ clknet_leaf_31_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5656__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _1948_ _2210_ _2226_ _1671_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7189_ _0012_ clknet_leaf_66_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5408__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6616__I _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7356__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4580__B _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3975__I _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6384__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4072__S _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4395__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6136__A2 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__A3 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5498__I1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6611__A3 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A2 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3910_ _3445_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4890_ _1039_ _1050_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_83_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3841_ _3375_ _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3885__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5078__S _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__A4 _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3772_ _3306_ _3307_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6560_ _0585_ _2509_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5511_ _1554_ _1555_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6491_ _1183_ _2467_ _2500_ _1097_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6127__A2 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4138__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ _1316_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7229__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5373_ _1317_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7112_ _3065_ _3069_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _0281_ _0506_ _0524_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7043_ as2650.r123\[0\]\[5\] _3006_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ _0309_ _0329_ _0372_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__C _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4161__I1 as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4186_ _0388_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3664__A3 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _2807_ _2810_ _2687_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3795__I _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _1540_ _0391_ _2744_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__A3 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _1137_ _1636_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6689_ _2677_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4301__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4852__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6054__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__B2 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5801__B2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__A3 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6293__A1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4040_ _3353_ _3562_ _3573_ _3517_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__A2 _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6045__A1 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ as2650.addr_buff\[2\] _1551_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6140__S1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _1098_ _1106_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _1040_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4359__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6612_ _1503_ _1599_ _1882_ _2602_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3824_ _3359_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3755_ _3126_ _3289_ _3290_ _3129_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6543_ _2493_ _2548_ _2549_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3686_ _3219_ _3221_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6474_ as2650.psu\[1\] _2466_ _1097_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _0783_ as2650.r123_2\[0\]\[6\] _1475_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6520__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4531__A1 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _0430_ _0506_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_87_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5287_ _0986_ _1376_ _1379_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7026_ _2983_ _2995_ _2996_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4238_ _0440_ _3270_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6036__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6587__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5011__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6511__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4522__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6785__B _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7067__A3 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_39_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6275__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6027__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6578__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6804__I _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4053__A3 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__I _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6502__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ as2650.stack\[2\]\[2\] _1329_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4513__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6190_ _0967_ _1936_ _2208_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4994__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ as2650.stack\[3\]\[3\] _1277_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7058__A3 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6266__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5072_ _0969_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4023_ as2650.r123\[1\]\[3\] as2650.r123_2\[1\]\[3\] _3136_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7417__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _1988_ _1995_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4856_ _3212_ _0512_ _1025_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _3327_ _3334_ _3340_ _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4787_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6741__A2 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4752__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ _2516_ _0772_ _2533_ _1159_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3738_ as2650.ins_reg\[5\] _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_118_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _0846_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5065__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3669_ _3203_ _3204_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4504__A1 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _0671_ _0682_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6388_ _2400_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _1409_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7009_ _2968_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4409__I _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6009__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4283__A3 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5232__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6732__A2 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6496__A1 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3932__B _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5703__I _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6799__A2 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6420__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6971__A2 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4054__I _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _0893_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ _1727_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__B net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4989__I _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _3128_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__S _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4572_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7360_ _0183_ clknet_leaf_30_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ _2172_ _2307_ _1799_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7291_ _0114_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4003__B _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6242_ _2256_ _2257_ _2258_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__I _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ _2189_ _2190_ _2191_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _1269_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ _1221_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4006_ _3422_ _3475_ _3533_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6411__A1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5957_ _1884_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6962__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _1066_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4973__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3776__A2 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _3328_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4839_ _3180_ _0866_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ as2650.psu\[3\] _2467_ _1652_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5951__C _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5150__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5523__I _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6402__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4192__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_54_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__A1 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7262__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6641__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _1136_ _2687_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _1837_ _1838_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _2749_ _2748_ _2750_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5742_ _1736_ _1775_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3758__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5673_ _0823_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7412_ _0235_ clknet_leaf_22_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _3221_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7343_ _0166_ clknet_3_0_0_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5380__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _0448_ _0693_ _0743_ _0715_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7274_ _0097_ clknet_leaf_50_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3930__A2 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _0677_ _3219_ _0678_ _0645_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__7121__A2 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _2239_ _2240_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5343__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6880__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__A3 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6156_ _0960_ _0759_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ as2650.stack\[4\]\[3\] _1222_ _1256_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _1125_ _2059_ _2005_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _1207_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3997__A2 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6935__A2 _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _1011_ _1584_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5518__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6699__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3921__A2 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput21 net21 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4578__B _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput32 net32 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput43 net43 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5674__A2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3685__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4332__I _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4340_ _3563_ _0537_ _0542_ _3352_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7103__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4271_ as2650.r0\[6\] _3145_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6010_ _0824_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4935__C _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6614__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6912_ _2302_ _2893_ _1788_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6843_ _2635_ _2825_ _2827_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4951__B _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6917__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6774_ _1940_ _2091_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _3312_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5725_ _1566_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5656_ _1487_ _1697_ _1698_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4607_ _0600_ _0687_ _0688_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5353__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7326_ _0149_ clknet_leaf_6_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3903__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4538_ _0338_ _0652_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ _0080_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4469_ _3311_ _0638_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5656__A2 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6208_ _1662_ _2216_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7188_ _0011_ clknet_leaf_67_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _2074_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5408__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6605__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A2 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7097__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6439__A4 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__A2 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4327__I _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__A4 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4622__A3 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A1 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3840_ _3351_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3771_ _3201_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _1557_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6490_ as2650.overflow _2466_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4138__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5372_ _0838_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _1759_ _1715_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7088__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _0281_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6835__A1 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7042_ _0424_ _3005_ _3007_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4254_ _0359_ _0457_ _0428_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4185_ _0346_ _0329_ _0360_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5110__I1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4074__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5777__B _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6452__I _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _2807_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _2742_ _2743_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5574__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3969_ _3503_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ _1601_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _2605_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5639_ _1562_ _1610_ _1588_ _1607_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4700__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _0132_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7323__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6826__A1 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4301__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5531__I _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__I1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4065__A1 _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7003__A1 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4368__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5580__A4 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5441__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4056__A1 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _1948_ _1987_ _1671_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5597__B _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _0672_ _1108_ _0877_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3803__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6611_ _1587_ _1617_ _1685_ _1874_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4359__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3823_ _3356_ _3358_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_92_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__I3 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6542_ _2510_ _0453_ _1083_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3754_ as2650.r0\[0\] _3125_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_leaf_9_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _1064_ _0847_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3685_ _3161_ _3210_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5616__I _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7346__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4520__I _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _0770_ _1478_ _1484_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5355_ _1006_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4306_ _0399_ _0429_ _0434_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5286_ as2650.stack\[0\]\[10\] _1377_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7025_ net21 _2986_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6284__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4237_ _3270_ _0371_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5351__I _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A1 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4047__A1 _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4099_ _0281_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ net33 _2794_ _2362_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5547__A1 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5011__A3 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__I _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5710__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__A2 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5140_ _0945_ _1276_ _1280_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5071_ _1233_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4022_ _3144_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A2 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5777__A1 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ _1798_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4515__I _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _0641_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5529__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _3219_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3806_ _3133_ _3341_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5774__C _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4786_ as2650.pc\[6\] _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4201__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6525_ _1653_ _0365_ _2532_ _2516_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3737_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4250__I _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _3432_ _2467_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3668_ as2650.idx_ctrl\[0\] _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_118_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _1450_ _1470_ _1471_ _1473_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6387_ _0993_ _2399_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3599_ as2650.halted net10 _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5338_ as2650.r123\[3\]\[6\] _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5269_ _0950_ _1363_ _1368_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7008_ _2969_ _2981_ _2982_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A2 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4283__A4 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__B _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4440__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6732__A3 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5940__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4160__I _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4259__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5759__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__B2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7191__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6184__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5931__A1 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _0489_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5166__I _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6310_ _2307_ _2317_ _2325_ _1850_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7290_ _0113_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6241_ as2650.pc\[8\] _1185_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _2189_ _2190_ _0750_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ as2650.stack\[4\]\[10\] _1244_ _1266_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5054_ as2650.stack\[5\]\[2\] _0942_ _1217_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5998__A1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4005_ _3536_ _3537_ _3538_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_84_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5956_ _1939_ _1979_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _3419_ _3462_ _0404_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5785__B _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4973__A2 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5887_ _0819_ _1906_ _1911_ _1655_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4838_ _0830_ _0998_ _1003_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6175__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5922__A1 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5076__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6508_ _3326_ _0847_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__A2 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6439_ _1869_ _1047_ _2449_ _2450_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4489__A1 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5150__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__A1 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6635__I _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6402__A2 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4413__A1 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4104__B _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7407__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6469__A2 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7150__B _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6641__A2 _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _1837_ _1838_ _1839_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _0376_ _0362_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5741_ _1737_ _1738_ _1758_ _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ _3554_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7411_ _0234_ clknet_leaf_20_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _0806_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_102_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7342_ _0165_ clknet_3_2_0_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _0381_ _0694_ _0692_ _0742_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7273_ _0096_ clknet_leaf_50_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4485_ _3364_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6224_ _1209_ as2650.stack\[3\]\[7\] as2650.stack\[2\]\[7\] _2241_ _2162_ _2242_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6155_ _1224_ net9 net1 as2650.pc\[5\] _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4486__A4 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4891__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3694__A2 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _1259_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6086_ _2103_ _2105_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__I _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5037_ _1151_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4643__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6396__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6988_ _1613_ _2965_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5939_ _1639_ _1943_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4703__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__A1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6699__A2 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput11 net11 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5534__I _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net51 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4594__B _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6623__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__I0 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6387__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6033__C _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5444__I _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ _3133_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6311__A1 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6075__B1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _0975_ _1322_ _2855_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ net34 _2794_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6378__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__I0 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3848__B _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6773_ _2625_ _2759_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3985_ _3494_ _3322_ _3382_ _3519_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5619__I _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5724_ _1738_ _1319_ _1752_ _1756_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _3316_ _1609_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4606_ _0719_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5586_ _0850_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6550__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7325_ _0148_ clknet_leaf_4_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ _0657_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5354__I _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7256_ _0079_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6302__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _0660_ _0631_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6302__B2 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _0818_ _2223_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7187_ _0010_ clknet_leaf_0_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4399_ _3392_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6138_ _2146_ _2147_ _1779_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6605__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _2087_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3602__I _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4616__A1 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A2 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4219__I1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7252__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4919__A2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7097__A2 _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__B1 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4607__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3830__A2 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5032__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6979__B _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _0902_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5174__I _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ _3066_ _3067_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3897__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4322_ _0402_ _0502_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7088__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5099__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7041_ as2650.r123\[0\]\[4\] _3006_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4253_ _0397_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4846__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5902__I _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ _3386_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4161__I3 as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4518__I _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7275__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4074__A2 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6825_ _2808_ _2773_ _2809_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5023__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4253__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ _0336_ _0348_ _2685_ _2719_ _2720_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5574__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3968_ _3502_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ net30 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3899_ _3434_ _3419_ _3430_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6523__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _1682_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5569_ _0860_ _0916_ _0861_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3888__A2 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7079__A2 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7308_ _0131_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6826__A2 _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7239_ _0062_ clknet_leaf_42_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4837__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4428__I _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A2 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A2 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__I _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A2 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6514__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6817__A2 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7298__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4338__I _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4056__A2 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _0826_ _1109_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _3208_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3822_ _3144_ _3357_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6610_ _1034_ _2599_ _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6541_ _2494_ _0470_ _2547_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3753_ as2650.r123\[1\]\[0\] as2650.r123_2\[1\]\[0\] _3288_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4801__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6505__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ _1741_ _3484_ _2479_ _2482_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3684_ _3186_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ as2650.r123_2\[0\]\[5\] _1481_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5354_ _3261_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4305_ _0449_ _0506_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5285_ _0981_ _1376_ _1378_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7024_ _0585_ _2960_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4236_ as2650.holding_reg\[5\] _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5492__A1 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4295__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__B _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4098_ _3402_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _2605_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5547__A2 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6744__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6739_ _1788_ _2709_ _2726_ _1083_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6412__B _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4711__I _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4158__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5235__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5086__I1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6306__C _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3797__A1 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6735__A1 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4597__I0 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5717__I _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7160__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7160__B2 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3721__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4269__S _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5070_ as2650.stack\[5\]\[6\] _1232_ _1227_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5474__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4021_ as2650.r123\[0\]\[3\] as2650.r123\[2\]\[3\] as2650.r123_2\[0\]\[3\] as2650.r123_2\[2\]\[3\]
+ _3142_ _3495_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_96_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6974__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5777__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _1989_ _1987_ _1993_ _1994_ _1753_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_80_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _3213_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3805_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _3139_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4785_ _0962_ _0956_ _0963_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4201__A2 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3736_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6524_ _3335_ _0848_ _2531_ _1653_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3667_ as2650.idx_ctrl\[1\] _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_106_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7151__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5406_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6386_ _1246_ _2371_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3598_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5337_ _1408_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5362__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ as2650.stack\[0\]\[3\] _1364_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7007_ net44 _2970_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4219_ _0394_ _0423_ _3447_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5199_ _1137_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6193__I _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__B1 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6965__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3610__I _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4976__B1 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6717__A1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__B2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6732__A4 _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3951__A1 _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4259__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7336__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6708__A1 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4195__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ _0757_ _3193_ _0649_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5931__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__A1 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__B _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7133__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _2085_ _2090_ _2132_ _2254_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6171_ _0538_ _0473_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _1268_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5447__A1 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5053_ _1220_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4004_ _3203_ _3299_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5955_ _1429_ _1938_ _1967_ _1462_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4906_ _1063_ _1072_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5886_ _1525_ _0750_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4973__A3 _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4837_ _1004_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5357__I _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5922__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3933__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6507_ _1095_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3719_ _3254_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7124__A1 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ _3156_ _1043_ _1686_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7209__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4210__B _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5092__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3605__I _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6369_ _2266_ _2381_ _2382_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__C _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7359__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5989__A2 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4661__A2 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6938__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6938__B2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6402__A3 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5610__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6651__I _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4177__A1 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__I _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4346__I _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_63_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5601__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _1759_ _1035_ _1773_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_76_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5671_ _1704_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5177__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4081__I as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7410_ _0233_ clknet_leaf_20_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4622_ _0676_ _0271_ _3162_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_124_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7341_ _0164_ clknet_leaf_17_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4553_ _0377_ _0651_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7106__A1 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__I _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7272_ _0095_ clknet_3_5_0_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4484_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5668__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _1919_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6154_ as2650.pc\[6\] net2 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ as2650.stack\[4\]\[2\] _0942_ _1256_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6085_ _2103_ _2105_ _0624_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6093__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _1205_ _1160_ _1062_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4643__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__B2 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6987_ _3171_ _1015_ _1604_ _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5938_ _1040_ _1938_ _1959_ _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_107_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5869_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3906__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput12 net12 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5659__A1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput23 net23 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6320__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7181__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3685__A3 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5682__I1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3938__C _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5725__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4570__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3756__S0 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4873__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6075__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6075__B2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6910_ _2769_ _2888_ _2891_ _1821_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _0883_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6505__B _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4389__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _1540_ _1499_ _2758_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3984_ _3324_ _3423_ _3518_ _3380_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6224__C _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ _1588_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5889__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _0585_ _0690_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5585_ _1615_ _1625_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5353__A3 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6550__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7324_ _0147_ clknet_leaf_5_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4536_ _3504_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7255_ _0078_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4467_ _3317_ _0635_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _1136_ _0921_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4398_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7186_ _0009_ clknet_leaf_67_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4695__B _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6137_ _1664_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5370__I _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _2088_ _2045_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_93_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5813__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__A2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5019_ as2650.psu\[1\] _1172_ _1174_ as2650.psu\[3\] _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6415__B _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__I _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3830__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6044__C _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5032__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6780__A2 _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4791__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6060__B _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6532__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _3181_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ _0511_ _0522_ _0523_ _0402_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4252_ _3298_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7040_ _2999_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__A2 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4183_ _3388_ _0358_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6048__A1 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _2799_ _0469_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5023__A2 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6755_ _2712_ _0348_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3967_ _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5706_ _1739_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _2635_ _2673_ _2675_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ _3325_ _3432_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5637_ _1492_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6523__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4534__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _1597_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7307_ _0130_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4519_ _0698_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5499_ _1549_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6287__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7238_ _0061_ clknet_leaf_54_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4837__A2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4709__I as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7169_ _1709_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3613__I _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__I _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6211__B2 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6762__A2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A1 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A2 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ _0647_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3821_ as2650.r123\[0\]\[1\] as2650.r123\[2\]\[1\] as2650.r123_2\[0\]\[1\] as2650.r123_2\[2\]\[1\]
+ _3142_ _3136_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6540_ _1683_ _0467_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3752_ as2650.psl\[4\] _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6471_ _1436_ _2480_ _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3683_ _3218_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6505__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4516__A1 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _0754_ _1477_ _1483_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _1416_ _1418_ _1419_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6269__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ _0399_ _0434_ _0432_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4119__I1 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5284_ as2650.stack\[0\]\[9\] _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7242__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7023_ _2961_ _1141_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4235_ _0431_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5492__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4166_ _0367_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__C _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4097_ _0287_ _3561_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7392__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _1230_ _2637_ _2786_ _2608_ _2792_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6744__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _1162_ _1163_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6738_ _1605_ _2711_ _2725_ _1787_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _1842_ _2658_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5095__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3608__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4507__A1 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6680__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__B2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A2 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4746__A1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_17_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6499__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7265__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6829__I _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5171__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5733__I _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3721__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ as2650.r0\[2\] _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5971_ _1899_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6974__A2 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4985__A1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4922_ _1081_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _0648_ _3318_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6726__A2 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4812__I _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3804_ _3335_ as2650.r123_2\[1\]\[7\] _3338_ _3339_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4784_ as2650.stack\[6\]\[5\] _0957_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6523_ as2650.psu\[4\] _2469_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3735_ _3270_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _0844_ _1099_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_109_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3666_ _3195_ _3201_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7151__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__B _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3872__B _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _3449_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5162__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _0990_ _1886_ _2397_ _2398_ _1591_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3597_ _3128_ _3132_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5336_ as2650.r123\[3\]\[5\] _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ _0944_ _1363_ _1367_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6662__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7006_ _0725_ _2976_ _2980_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _1323_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4149_ as2650.r123\[2\]\[3\] _3451_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__B _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4976__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6717__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7288__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3951__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5553__I _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4900__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__I _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6653__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3801__I _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5208__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6956__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__I _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7148__C _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5891__C _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6341__B1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6170_ _2141_ _2143_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5121_ as2650.stack\[4\]\[9\] _1241_ _1266_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3912__S _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6644__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5447__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ as2650.stack\[5\]\[1\] _1219_ _1217_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4807__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ _3437_ _3361_ _3503_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_133_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3711__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4905_ _1073_ _1071_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5885_ _1433_ _1909_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3630__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__I _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4836_ _3364_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5383__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6506_ _0334_ _1665_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3933__A2 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3718_ _3253_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4698_ _3262_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6437_ _3202_ _3310_ _1008_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3649_ _3184_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5373__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6883__A1 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6368_ as2650.addr_buff\[3\] _0624_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ _0980_ _1397_ _1399_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6299_ _1528_ _2281_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6418__B _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6938__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7060__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3621__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4177__A2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3924__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__I _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6323__B1 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6874__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5677__A2 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__B _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6929__A2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3860__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7051__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3612__A1 _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _1711_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4621_ _3192_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5365__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _0163_ clknet_leaf_30_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _0290_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__C _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7271_ _0094_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4483_ _3182_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5668__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6865__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _2199_ as2650.stack\[1\]\[7\] as2650.stack\[0\]\[7\] _1252_ _2240_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4340__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6153_ _1896_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5921__I _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _1258_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6084_ net9 _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _1152_ _1155_ _1203_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5840__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7042__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _1820_ _1415_ _1143_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5937_ _0900_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _3247_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4819_ as2650.stack\[6\]\[11\] _0983_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5799_ _1324_ _1820_ _1821_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7326__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput13 net49 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6856__A1 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6927__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4331__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6084__A2 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4447__I _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5831__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7033__A1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5347__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4910__I _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5898__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__A2 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4322__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3756__S1 _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4357__I _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6075__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4086__A1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _1232_ _2637_ _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2268_ _2741_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3983_ _3353_ _3504_ _3516_ _3517_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _1696_ _1754_ _0851_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ _0869_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7349__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4604_ _0785_ _0691_ _0789_ _0698_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5889__A2 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4010__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5584_ _1445_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7323_ _0146_ clknet_leaf_5_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4535_ as2650.r0\[3\] _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6838__B2 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7254_ _0077_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4466_ _3348_ _0639_ _0658_ _0634_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ _1548_ _1908_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4313__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7185_ _0008_ clknet_leaf_0_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5651__I _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _0389_ _0579_ _0581_ _3388_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_86_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _2009_ _2151_ _2154_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4267__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ as2650.pc\[3\] net8 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4077__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5018_ as2650.psu\[4\] _1184_ _1187_ net27 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4616__A3 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__A3 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _2908_ _2944_ _2947_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4730__I _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A2 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4068__A1 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A1 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4640__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4320_ _0419_ _0504_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7172__B _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4251_ _0454_ _0373_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4182_ _0363_ _3322_ _0364_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__A1 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6823_ _2799_ _0469_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5023__A3 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ _2739_ _2740_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3966_ _3497_ _3500_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _1511_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ net29 _2674_ _2362_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3897_ _3414_ _3418_ as2650.psl\[3\] _3432_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5636_ _1650_ _1668_ _1681_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4534__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ _1599_ _1608_ _1611_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7306_ _0129_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4518_ _0664_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5498_ _1324_ _1548_ _1523_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6287__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _0060_ clknet_leaf_43_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ _3159_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5381__I _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7168_ _1313_ _3105_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6119_ _1945_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7099_ _2471_ _2462_ _3057_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5556__I _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5789__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__B _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7194__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4461__A1 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6850__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ _3126_ _3354_ _3355_ _3130_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7167__B _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3751_ _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__I _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _1855_ _3492_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3682_ as2650.ins_reg\[7\] _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5421_ as2650.r123_2\[0\]\[4\] _1481_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4516__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ _1420_ _0623_ _0917_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5283_ _1361_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7022_ _2983_ _2992_ _2993_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4234_ _0400_ _0407_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4165_ _3127_ _0368_ _0369_ _3131_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4096_ _0294_ _0297_ _0300_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6441__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4452__A1 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6806_ _1900_ _2136_ _2791_ _2250_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4998_ _3372_ _3438_ _0530_ _1164_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5547__A4 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6737_ _2718_ _2724_ _2659_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3949_ _3456_ _3483_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5952__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6668_ _0317_ _1488_ _1489_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5619_ _1046_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6599_ _0980_ _2591_ _2593_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3624__I as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6000__I _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6680__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A2 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4746__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5943__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4190__I _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5171__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_57_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3721__A3 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6120__A1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6959__B1 _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__I _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6423__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5970_ _1990_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _1077_ _1079_ _1084_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_79_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4985__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _0914_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6726__A3 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3803_ _3139_ as2650.r123\[1\]\[7\] _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4783_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5196__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _0751_ _0423_ _2457_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3734_ _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6453_ _1114_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3665_ _3196_ _3200_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5924__I _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__C _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _0895_ _1449_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6384_ _1888_ _2373_ _1889_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3596_ _3131_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5335_ _1407_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5266_ as2650.stack\[0\]\[2\] _1364_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6111__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7005_ _2972_ _0741_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4217_ _0395_ _0401_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_102_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5197_ _1025_ _1304_ _1312_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4673__A1 as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4148_ _3447_ _0307_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_95_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6414__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ _3584_ _0263_ _0266_ _0273_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4425__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4208__C _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6178__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__C _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5925__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6350__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__B2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__A3 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4664__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4118__C _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4913__I _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6169__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5392__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6341__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__B2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5120_ _1267_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6575__I _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5051_ _0936_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A1 _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4002_ _3423_ _3510_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4095__I _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _1969_ _1970_ _1976_ _1927_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4823__I _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _0559_ _0564_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5884_ _1907_ _1908_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3630__A2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _0835_ _0903_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5907__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4766_ as2650.pc\[3\] _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3717_ _3179_ _3160_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6505_ _1741_ _0307_ _2479_ _2513_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7485_ net47 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _0867_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5654__I _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7074__C _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6332__A1 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5135__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3648_ _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6436_ _1055_ _1058_ _2447_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6883__A2 _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _1131_ _1739_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4894__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5318_ as2650.stack\[1\]\[9\] _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6298_ _0869_ _2309_ _2311_ _2220_ _2313_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_102_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5438__A3 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ as2650.r123_2\[1\]\[4\] _1354_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3902__I _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_2_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6399__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7255__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4949__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5829__I _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3621__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6571__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A2 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6323__B2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6874__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4885__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5513__B _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6328__C _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6344__B _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5365__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6562__A1 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4551_ _0362_ _0709_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7270_ _0093_ clknet_leaf_50_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4482_ _3209_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5407__C _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6314__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _1457_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6865__A2 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3679__A2 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _0964_ _2170_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ as2650.stack\[4\]\[1\] _1219_ _1256_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4818__I _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _3140_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3722__I _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4628__A1 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5034_ _1093_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7278__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7042__A2 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6985_ _3317_ _2960_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _3506_ _1511_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _1616_ _1630_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4818_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6553__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5798_ _1825_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4749_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5384__I _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6305__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6305__B2 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net14 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput25 net25 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5659__A3 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6419_ _0824_ _2428_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xoutput36 net36 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7399_ _0222_ clknet_leaf_36_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4867__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6429__B _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3632__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A3 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3842__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7033__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5347__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__I _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7426__D _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4570__A3 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4858__A1 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7420__CLK clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__I _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4086__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6083__I0 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5035__B2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6770_ _1857_ _2738_ _2741_ _2693_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3982_ _3168_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3597__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5721_ _1093_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5652_ _1689_ _1693_ _1694_ _1695_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6535__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4603_ _0715_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5583_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4010__A2 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7322_ _0145_ clknet_leaf_2_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4534_ _0686_ _0723_ _0724_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6838__A2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7253_ _0076_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4465_ _3510_ _0644_ _0654_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6204_ _1234_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7184_ _0007_ clknet_leaf_6_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4396_ _3344_ _3550_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5510__A2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6135_ _0871_ _1945_ _1946_ _3233_ _1105_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ as2650.pc\[3\] _0335_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4077__A2 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__A2 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6968_ _1542_ _2945_ _2946_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6774__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5577__A2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4216__C _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5919_ _0868_ _1937_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6899_ _0975_ _2700_ _2881_ _2699_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4458__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__B _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5265__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3815__A2 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4240__A2 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7009__I _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4250_ _3543_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ _3257_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4059__A2 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5199__I _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6822_ _1187_ _0548_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7316__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5559__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5023__A4 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6753_ _2707_ _2710_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3965_ _3126_ _3498_ _3499_ _3130_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5704_ _1295_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6508__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6684_ _2605_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3896_ as2650.carry _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5635_ _1647_ _1651_ _1667_ _1680_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_136_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5566_ _1494_ _1612_ _3212_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3742__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7305_ _0128_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4517_ _0686_ _0706_ _0708_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5497_ _0316_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5662__I _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7236_ _0059_ clknet_leaf_42_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4448_ _0640_ _3252_ _3401_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5495__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4278__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7167_ _1313_ _1643_ _3102_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4379_ _3343_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_98_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _1988_ _2137_ _1996_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _2465_ _0773_ _3056_ _2471_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6049_ as2650.stack\[6\]\[3\] _1921_ _1969_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_73_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__S _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4470__A2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6747__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4222__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4741__I _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3981__A1 _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7172__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4289__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6986__A1 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6336__C _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6738__A1 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__B _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4213__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3750_ _3134_ _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6071__C _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7163__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3681_ _3172_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _0737_ _1477_ _1482_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6910__A1 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5351_ _0316_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__I _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4302_ _0502_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5282_ _1362_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4119__I3 as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7021_ net20 _2986_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4233_ _0398_ _0418_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4164_ as2650.r0\[5\] _3143_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5229__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6527__B _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__I as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4095_ _3480_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3730__I _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6977__B2 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__C _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout52_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__A3 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6729__A1 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6805_ _1230_ _2787_ _2789_ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__I _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4997_ _1165_ _0799_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4561__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _1131_ _2653_ _2723_ _1492_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3948_ _3482_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7154__A1 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _2649_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3879_ _3268_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5618_ _1297_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6901__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6901__B2 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ as2650.stack\[7\]\[9\] _2592_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__I _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5549_ _0851_ _1055_ _1555_ _3165_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7219_ _0042_ clknet_leaf_59_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6172__B _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3954__A1 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7145__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__3721__A4 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6959__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5631__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4920_ _1063_ _1085_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _3273_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6726__A4 _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3802_ _3128_ _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4782_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3945__A1 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _2493_ _2527_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7136__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3733_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _1046_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3664_ as2650.cycle\[6\] _3154_ _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_118_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5698__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _1463_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3595_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3725__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6383_ _1800_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4370__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6101__I _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ as2650.r123\[3\]\[4\] _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5265_ _0939_ _1363_ _1366_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _2969_ _2978_ _2979_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4216_ _0402_ _0398_ _0413_ _0420_ _3400_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ _1109_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4673__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5870__A1 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4147_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4078_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5622__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4492__S _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5925__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3936__A1 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ net31 _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7184__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6011__I _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6638__B1 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4113__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__A3 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4664__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__S _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4416__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5613__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7429__D _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__B1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6122__S _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _1218_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4104__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _3534_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5852__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4655__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _1971_ _1973_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6524__C _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _1064_ _0558_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5883_ _1510_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4834_ _0622_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5000__I as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7109__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _0945_ _0933_ _0946_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6580__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6504_ _2510_ _2511_ _2512_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3716_ _3210_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4591__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7484_ net47 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4696_ _0870_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6435_ _1063_ _2445_ _2446_ _1501_ _1613_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3647_ as2650.ins_reg\[4\] _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6332__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _2378_ _2372_ _0832_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _1382_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6297_ _0979_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6096__A1 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5603__C _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _0737_ _1350_ _1355_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4286__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5843__A1 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _3199_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3909__A1 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4582__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6323__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4885__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6676__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5513__C _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4924__I _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6344__C _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5755__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5365__A3 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6562__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4550_ _0686_ _0737_ _0739_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _0639_ _0625_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6220_ as2650.stack\[7\]\[7\] as2650.stack\[4\]\[7\] as2650.stack\[5\]\[7\] as2650.stack\[6\]\[7\]
+ _0928_ _2237_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3679__A3 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__A2 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6151_ _1229_ _2130_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _1257_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ _2063_ _2101_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5825__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5033_ _1157_ _1159_ _1201_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_111_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6984_ _2961_ _2462_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6250__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5935_ _1955_ _1957_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _0889_ _1432_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5797_ _1548_ _1820_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6553__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5665__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4564__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4679_ _0849_ _0852_ _0856_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4316__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ _2288_ _2429_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput15 net15 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput26 net26 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ _0221_ clknet_leaf_35_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput37 net37 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4867__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6349_ _0987_ _1936_ _2363_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3913__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7222__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5816__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7372__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6241__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6792__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__C _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__A1 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6355__B _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__I _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6083__I1 as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3981_ _3507_ _3509_ _3376_ _3515_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__S _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ _1753_ _1663_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3597__A2 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5651_ _1472_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6535__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _0587_ _0758_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5582_ _0537_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7321_ _0144_ clknet_leaf_3_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4533_ as2650.r123_2\[2\]\[2\] _0707_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__A1 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _0075_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7245__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6203_ _0965_ _2148_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4829__I _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7183_ _0006_ clknet_leaf_7_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3733__I _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4395_ _0585_ _0314_ _0364_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _1433_ _2152_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6471__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5016_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5026__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _1542_ _2929_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6774__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4785__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5918_ _0936_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6898_ _1664_ _2265_ _2880_ _1672_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5849_ _0843_ _0846_ _3246_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5395__I _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__A2 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5888__I1 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3643__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7115__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5265__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6462__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6175__B _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4474__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5519__B _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _3324_ _0365_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6085__B _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4384__I _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6205__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6821_ _1126_ _2641_ _2617_ _2805_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6813__B _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ net32 _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3964_ as2650.r0\[2\] _3331_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5703_ _1570_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6683_ _1219_ _2637_ _2672_ _2608_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3895_ _3410_ _3420_ _3427_ _3430_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3728__I _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6508__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5634_ _1310_ _1678_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3990__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5565_ _0317_ as2650.addr_buff\[7\] _3307_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7304_ _0127_ clknet_leaf_53_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3742__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4516_ as2650.r123_2\[2\]\[1\] _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5496_ _1546_ _1526_ _1547_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7235_ _0058_ clknet_leaf_43_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4447_ _3161_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6692__A1 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _3083_ _3116_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4378_ _0464_ _0529_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _1903_ _2131_ _2136_ _1900_ _2048_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_115_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _1698_ _3055_ _2465_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6444__A1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _2023_ _2068_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7257__D _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7172__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5183__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5183__B2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4930__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__B2 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6684__I _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6435__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6435__B2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5789__A3 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6986__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4997__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6738__A2 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4932__I _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6352__C _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ _3178_ _3193_ _3206_ _3215_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7163__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5763__I _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6910__A2 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4921__A1 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5350_ _1107_ _1298_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ as2650.holding_reg\[6\] _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ _1375_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _1728_ _2960_ _2991_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _0433_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4163_ as2650.r123\[1\]\[5\] as2650.r123_2\[1\]\[5\] _3495_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6426__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4094_ _0271_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6977__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7433__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__A2 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6804_ _1443_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4996_ _3211_ _3587_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6735_ _2653_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3947_ _3474_ _3477_ _3481_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6666_ _1173_ _2613_ _2655_ _1826_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3878_ _3253_ _3295_ _3411_ _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_104_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5617_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6597_ _2576_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5673__I _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6901__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3715__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ _3232_ _0409_ _1024_ _1029_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_118_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5479_ as2650.addr_buff\[2\] _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7218_ _0041_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5622__B net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7149_ _3095_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5114__S _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6417__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6417__B2 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7090__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5848__I _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout50 net36 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7145__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5583__I _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__B _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4903__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3706__A2 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5459__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4927__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3831__I _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6408__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6959__A2 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5631__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4662__I _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4850_ _1012_ _1015_ _1016_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3801_ _3336_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _1856_ _0391_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3732_ as2650.ins_reg\[3\] as2650.ins_reg\[2\] _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _1145_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3663_ _3197_ _3198_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6895__A1 _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6382_ _2370_ _2374_ _2379_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3594_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _1406_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5264_ as2650.stack\[0\]\[1\] _1364_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6538__B _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7003_ net43 _2970_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4215_ _3579_ _0416_ _0418_ _0419_ _3403_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _1321_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5870__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4146_ _3521_ _0313_ _0351_ _3283_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3881__A1 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7072__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4077_ as2650.holding_reg\[3\] _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3897__B as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6718_ _2676_ _2678_ _2697_ _2706_ _1591_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3936__A2 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ net52 net28 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7329__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6886__A1 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6638__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6638__B2 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4113__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5310__A1 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7063__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6810__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5613__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A1 _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6911__B _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5377__B2 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6630__C _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5527__B _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3826__I _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6877__A1 _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6202__I _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4352__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6629__A1 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4104__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6077__C _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4000_ _3533_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5852__A2 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3863__A1 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__S _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7054__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _0893_ as2650.stack\[3\]\[1\] as2650.stack\[2\]\[1\] _1974_ _1467_ _1975_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_111_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5488__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _0514_ _1065_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5882_ _3373_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _3194_ _0757_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6821__B _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4764_ as2650.stack\[6\]\[2\] _0934_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7109__A2 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6503_ _1827_ _0349_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3715_ _3187_ _3249_ _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7483_ net47 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3736__I _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4695_ as2650.psu\[5\] _0873_ _0875_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6868__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6868__B2 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _1025_ _3266_ _0655_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3646_ as2650.ins_reg\[2\] _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5540__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _1900_ _2378_ _2373_ _1903_ _1462_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5316_ _1383_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _0974_ _0969_ _2221_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__B _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6096__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ as2650.r123_2\[1\]\[3\] _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5843__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5178_ _1305_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3854__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4129_ net8 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6020__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__A1 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__A3 _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3646__I as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5861__I _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6178__B _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__I _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A1 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5834__A2 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5598__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5365__A4 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5770__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7028__I _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4480_ _0671_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3679__A4 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6150_ _0962_ _1983_ _2169_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6088__B _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5101_ as2650.stack\[4\]\[0\] _1208_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__I _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6081_ _0335_ _2061_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5125__I1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _1121_ _0587_ _1115_ _1158_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7027__A1 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _2959_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6250__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _1955_ _1957_ _1558_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4261__A1 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5865_ _0890_ _1888_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4816_ as2650.pc\[11\] _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5796_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4013__A1 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4564__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _0895_ _0899_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4678_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6417_ _2119_ as2650.stack\[3\]\[12\] as2650.stack\[2\]\[12\] _1929_ _1468_ _2430_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_123_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4316__A2 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3629_ _3161_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5513__A1 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _0220_ clknet_leaf_35_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput16 net16 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ _2129_ _2361_ _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__I1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6279_ _2250_ _2294_ _2295_ _2252_ _1981_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4246__B _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6241__A2 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6792__A3 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6461__B _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4760__I _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5752__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6687__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5805__B _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4307__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__I1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7197__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6480__A2 _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6355__C _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ _3509_ _3514_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A1 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5766__I _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _3297_ _1689_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _0589_ _0651_ _0758_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5743__A1 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _0381_ _0488_ _0591_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_129_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _0143_ clknet_leaf_67_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _0278_ _0722_ _0667_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7251_ _0074_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6597__I _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4463_ _0655_ _3166_ _0629_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6202_ _1893_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7182_ _0005_ clknet_leaf_6_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4394_ _3380_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _0832_ _2131_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _0953_ net9 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ net2 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A3 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _1538_ _2646_ _2928_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5917_ _0887_ as2650.ins_reg\[2\] _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4785__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__A1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ _1525_ _0751_ _2879_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _1594_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5779_ _1810_ _1053_ _1802_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6175__C _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5586__I _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5519__C _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6150__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _2641_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _2086_ _2737_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3963_ as2650.r123\[1\]\[2\] as2650.r123_2\[1\]\[2\] _3136_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _1736_ _1038_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6682_ _1084_ _2664_ _2671_ _1094_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3894_ _3429_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _0909_ _1676_ _1083_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5564_ _1440_ _1609_ _1610_ _0918_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_129_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4515_ _0684_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7303_ _0126_ clknet_leaf_44_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3742__A3 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5495_ _3234_ _1523_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ _0636_ _0637_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6141__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7234_ _0057_ clknet_leaf_42_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6141__B2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6692__A2 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7165_ as2650.psu\[2\] _3113_ _3115_ _3096_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4377_ _0556_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6116_ _2133_ _2135_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7096_ _1128_ _2018_ _0804_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6047_ as2650.stack\[7\]\[3\] _1922_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4455__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5955__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _2389_ _2905_ _2906_ _2907_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__3805__I1 as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__B2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5183__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6380__B2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4930__A2 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A1 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6683__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4485__I _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7235__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4300_ _0480_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6123__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ _0977_ as2650.stack\[0\]\[8\] _1362_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ _0399_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4685__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4162_ _3336_ _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6426__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4093_ as2650.holding_reg\[3\] _3254_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_83_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4437__A1 _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6803_ _2139_ _2783_ _2788_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ _3132_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _0337_ _0349_ _2721_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3946_ _3478_ _3480_ _3461_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ _2650_ _2651_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3877_ _3291_ _3293_ _3412_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_137_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4998__C _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _0810_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6362__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6596_ _2577_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5547_ _3260_ _1032_ _0902_ _1491_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__3715__A3 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5478_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4429_ _3277_ _3226_ _3224_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7217_ _0040_ clknet_leaf_55_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4676__A1 _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6718__C _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7148_ _3096_ _3098_ _3101_ _2736_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7079_ _0560_ _1701_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7090__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5928__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout51 net33 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__I _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6353__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6353__B2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4903__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3706__A3 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4667__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6408__A2 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7081__A2 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4943__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5919__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ as2650.ins_reg\[0\] _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4780_ as2650.pc\[5\] _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ _3205_ _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_35_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3662_ as2650.cycle\[0\] _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5147__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6344__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _3438_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5401_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6895__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _1319_ _2388_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3593_ as2650.ins_reg\[0\] _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5332_ as2650.r123\[3\]\[3\] _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5263_ _0892_ _1363_ _1365_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4658__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7002_ _1713_ _2976_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4214_ _0301_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5194_ _1320_ _0873_ _1311_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7400__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4145_ _3313_ _0345_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5014__I _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3881__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7072__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4076_ _3556_ _3559_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3897__C _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6273__C _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4830__A1 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6583__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5386__A2 as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ net10 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6717_ _0942_ _2698_ _2704_ _1800_ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3929_ _3459_ _3461_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6648_ _1787_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5138__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6335__A1 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6886__A2 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6579_ _0938_ _2578_ _2581_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5633__B _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5125__S _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6448__C _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4113__A3 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7063__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4763__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5377__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7118__A3 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__A1 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4938__I _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__A3 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6374__B _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__I _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5950_ _1456_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _1064_ _0559_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5881_ _0833_ _1898_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4832_ _1000_ _1001_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6565__A1 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4763_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4040__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _1683_ _0313_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6317__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3714_ _3190_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7482_ net46 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4694_ _0873_ _0876_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _1080_ _1006_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3645_ _3180_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6364_ _2375_ _2377_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5540__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5315_ _1396_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6295_ _1960_ _2310_ _1441_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5246_ _1347_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5843__A3 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5177_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4128_ _0289_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5679__I _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ as2650.holding_reg\[2\] _3415_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6005__B1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5628__B _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__A1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4319__B1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6859__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4334__A3 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7036__A2 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__I _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__A1 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5598__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6547__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3837__I _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4022__A2 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5070__I1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5770__A2 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4668__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6088__C _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6080_ _0335_ _2061_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5031_ _1053_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7027__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7319__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _1171_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_50_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _1885_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6538__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5448__B _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4815_ _0987_ _0982_ _0988_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5795_ _1747_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4746_ _0920_ _0926_ _0929_ _3264_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__3772__A1 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4677_ _0857_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6416_ _1212_ as2650.stack\[1\]\[12\] as2650.stack\[0\]\[12\] _2072_ _2429_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3628_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5513__A2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6710__A1 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _0219_ clknet_leaf_36_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput17 net17 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_115_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6347_ _0883_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _2172_ _2263_ _2180_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5277__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ _0981_ _1341_ _1343_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6777__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__B2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6529__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7129__I _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5052__I1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__I _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _0591_ _0652_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5743__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ _3514_ _3567_ _0334_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3754__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4531_ _3545_ _0709_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7250_ _0073_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ _3157_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6201_ _1896_ _2217_ _2218_ _2180_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7181_ _0004_ clknet_leaf_7_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4393_ _3517_ _0586_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6132_ _1948_ _2136_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6827__B _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _0375_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6759__A1 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7291__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6965_ net40 _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5431__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__I _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4861__I _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ _1442_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _2667_ _2875_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5982__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _0675_ _0821_ _0862_ _1834_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6931__A1 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5778_ _3229_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4729_ _3185_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5692__I _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7379_ _0202_ clknet_leaf_15_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4101__I _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__B _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__I _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6998__A1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__B _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6472__B _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4225__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7175__A1 as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7175__B2 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5186__B1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__B _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6989__A1 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5978__S _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5661__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4216__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _2087_ _2708_ _2088_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ _3144_ _3496_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ _1735_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7166__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6681_ _1219_ _2665_ _2670_ _2623_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3893_ _3218_ _3428_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5632_ _1143_ _1642_ _1674_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__6913__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3727__A1 _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__B _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5563_ _1048_ _1035_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7302_ _0125_ clknet_leaf_44_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6401__I _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ _3484_ _0627_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5494_ _1187_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7233_ _0056_ clknet_leaf_56_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4445_ _0629_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4152__A1 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7164_ _3066_ _3114_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4376_ _0458_ _0529_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6557__B _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__B _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _2085_ _2090_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3760__I _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7095_ _0577_ _3038_ _1204_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _2024_ as2650.stack\[5\]\[3\] as2650.stack\[4\]\[3\] _2025_ _2068_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5888__S _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__A2 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _2908_ _2905_ _2907_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_74_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5955__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3966__A1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _2858_ _2860_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6904__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__A2 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4391__A1 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__A3 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6132__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4766__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7142__I _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4446__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5643__A1 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6981__I _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A3 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6199__A2 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7148__A1 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__I _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4134__A1 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4230_ _0414_ _0295_ _0398_ _0303_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4685__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ as2650.r123\[0\]\[5\] as2650.r123\[2\]\[5\] as2650.r123_2\[0\]\[5\] as2650.r123_2\[2\]\[5\]
+ _3143_ _3495_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4092_ _3254_ _0288_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4437__A2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _0872_ _1768_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4994_ _0539_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5937__A2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6733_ _2685_ _2719_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3945_ _3479_ _3218_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6664_ _2650_ _2651_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3876_ as2650.holding_reg\[0\] _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5615_ _1655_ _1656_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4360__B _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6362__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7374__D _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6595_ _2590_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5546_ _3308_ _1496_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _1532_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4125__A1 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7216_ _0039_ clknet_leaf_9_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4428_ _3197_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4586__I _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7147_ _3099_ _3100_ net27 _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _0560_ _3344_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7078_ _1700_ _0567_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ _0941_ _2010_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_5_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net29 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4667__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7202__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_90 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_127_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _3146_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3661_ _3152_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6344__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4355__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _1465_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6380_ _1761_ _2392_ _2393_ _2006_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3592_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5331_ _1405_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5790__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5262_ as2650.stack\[0\]\[0\] _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7001_ _2972_ _0726_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4213_ _3270_ _0327_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5193_ _1319_ _1303_ _0447_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3961__S0 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4144_ _3392_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4075_ _0270_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6280__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__C _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout50_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6032__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _1092_ _1147_ _1062_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5965__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6716_ _2677_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4594__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3928_ _3408_ _3433_ _3462_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ _2636_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3859_ _3315_ _3384_ _3394_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6335__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6578_ as2650.stack\[7\]\[1\] _2579_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5529_ _3173_ _3279_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6099__B2 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4649__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5846__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5205__I _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4113__A4 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5875__I _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4954__I _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7054__A3 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _1069_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _0888_ _1432_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _0844_ _0800_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4762_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6501_ _1425_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3713_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7481_ net46 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6317__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4328__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ _1437_ _2443_ _3304_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3644_ _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7248__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4879__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6363_ _2333_ _2336_ _2376_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5314_ _1237_ as2650.stack\[1\]\[8\] _1383_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6294_ _1529_ _2268_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _0723_ _1350_ _1353_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _0903_ _1033_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4864__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4127_ _0331_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6253__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4058_ _3415_ _3502_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_80_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6556__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4567__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4319__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3943__I _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4774__I _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4558__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A3 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ _0822_ _1198_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4684__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _3238_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6786__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5932_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _3138_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4797__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4261__A3 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5863_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4814_ as2650.stack\[6\]\[10\] _0983_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5794_ _1748_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5210__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4676_ _3134_ _0812_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6415_ _2288_ _2426_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3627_ as2650.ins_reg\[5\] _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7395_ _0218_ clknet_leaf_35_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6710__A2 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6279__C _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net52 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6346_ _2331_ _2339_ _2360_ _2206_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _2263_ _2283_ _2293_ _1850_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__A1 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ as2650.stack\[2\]\[9\] _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5911__C _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6295__B _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5159_ as2650.stack\[3\]\[10\] _1290_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5029__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7413__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__A2 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5752__A3 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4769__I _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5268__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A1 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__A1 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4779__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_91_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _0689_ _0718_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3754__A2 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4951__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4461_ _3370_ _0651_ _0643_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6200_ _1903_ _2210_ _2048_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7180_ _0003_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4392_ _3572_ _0587_ _0593_ _3168_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _2148_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6062_ _1225_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5013_ as2650.psu\[2\] _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6208__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7436__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6964_ net39 _2925_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5431__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1887_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6895_ _2855_ _2856_ _1084_ _2877_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4363__B _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3993__A2 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5846_ _1417_ _1867_ _1868_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5777_ _3228_ _0825_ _1413_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4728_ _0857_ _0900_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4942__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5906__C _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _3337_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7378_ _0201_ clknet_leaf_15_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6329_ _0979_ _2312_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__A1 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3984__A2 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4499__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6135__B1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6686__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6438__A1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6989__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6610__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3961_ as2650.r123\[0\]\[2\] as2650.r123\[2\]\[2\] as2650.r123_2\[0\]\[2\] as2650.r123_2\[2\]\[2\]
+ _3142_ _3495_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5700_ _1149_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _2666_ _1951_ _2669_ _2626_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3892_ _3186_ as2650.ins_reg\[6\] _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5631_ _1412_ _1584_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _1502_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__C _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7301_ _0124_ clknet_leaf_44_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4513_ _0626_ _0702_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5493_ _1544_ _1526_ _1545_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7232_ _0055_ clknet_leaf_59_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4444_ _3166_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7163_ _1130_ _3105_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4152__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4375_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6114_ _1224_ _0377_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5461__C _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7094_ _0528_ _3036_ _1085_ _3038_ _3052_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _1869_ _2058_ _2066_ _2008_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3663__A1 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _1494_ _2390_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7157__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _2274_ _2858_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5168__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6365__B1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6117__B1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6668__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__A4 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__A3 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A2 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6840__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4446__A3 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5643__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__I _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4782__I _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7148__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4731__B _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5118__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6659__A1 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7281__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4957__I _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4134__A2 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3861__I _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5054__S _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ _3562_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7084__A1 _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _3579_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4692__I _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _2628_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _0588_ _0567_ _3361_ _3506_ _0330_ _0377_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_90_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6732_ _1532_ _3547_ _3549_ _3551_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3944_ _3249_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6663_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3875_ _3407_ _3253_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6898__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5614_ _1509_ _1657_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__6898__B2 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _1237_ as2650.stack\[7\]\[8\] _2577_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5545_ _3175_ _1590_ _1592_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5570__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5476_ _3568_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ _0605_ _0615_ _0620_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7215_ _0038_ clknet_leaf_9_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3771__I _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ _3095_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4676__A3 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A2 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4358_ as2650.holding_reg\[7\] _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4088__B _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3884__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7075__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6122__I0 as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7077_ _0501_ _1701_ _3035_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _3572_ _0481_ _0492_ _3323_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6822__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _1988_ _2049_ _1996_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__A1 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4107__I _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4061__A1 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout53 net26 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6338__B1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6478__B _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5382__B _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4777__I _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5313__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__A1 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6992__I _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__A1 _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3627__A1 as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5401__I _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_80 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_91 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4052__A1 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__B _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5049__S _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6232__I _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ as2650.cycle\[5\] as2650.cycle\[4\] _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4355__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3591_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ as2650.r123\[3\]\[2\] _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4687__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _1361_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7000_ _2959_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4212_ as2650.holding_reg\[4\] _3415_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5192_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7057__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4143_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3961__S1 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ _3287_ _0279_ _0280_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6280__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7177__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4291__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6568__B1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__A1 _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4976_ _1094_ _1140_ _1142_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6570__C _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ _0943_ _2700_ _2703_ _2699_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4371__B _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3927_ _3459_ _3461_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6142__I _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ _1554_ _1579_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3858_ _3391_ _3393_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _0891_ _2578_ _2580_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3789_ as2650.psl\[3\] _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5528_ _3479_ _1574_ _1576_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5459_ _0999_ _1417_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5846__A2 _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7048__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__B _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ _1696_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3609__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3676__I _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4300__I _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3848__A1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_2_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__I _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4830_ _3436_ _0645_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4025__A1 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5773__A1 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3712_ as2650.ins_reg\[6\] _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6500_ _2454_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7480_ net46 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _0802_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3643_ as2650.ins_reg\[3\] _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6431_ _3236_ _3240_ _3281_ _3276_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5525__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4328__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ as2650.pc\[10\] _0539_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4879__A3 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5313_ _0971_ _1390_ _1395_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6293_ _2053_ _2299_ _2308_ _0818_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ as2650.r123_2\[1\]\[2\] _1351_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _1128_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _3422_ _3475_ _3511_ _3534_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_111_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _3584_ _0263_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4264__A1 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5041__I _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6005__A2 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4880__I _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4016__A1 _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4567__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _0711_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ _2458_ _2615_ _2619_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__C _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5119__I1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6492__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6475__C _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4255__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4007__A1 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__I0 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5507__A1 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4030__I _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4965__I _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6385__C _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6980_ _2957_ _2958_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4246__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6786__A3 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _3371_ _1913_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5796__I _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _1048_ _1645_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4813_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5793_ _1822_ _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4744_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4675_ _0858_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7365__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3626_ as2650.ins_reg\[4\] as2650.ins_reg\[6\] as2650.ins_reg\[7\] _3162_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6414_ as2650.stack\[7\]\[12\] _1455_ _1974_ as2650.stack\[6\]\[12\] _1968_ _2427_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6171__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7394_ _0217_ clknet_leaf_52_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput19 net19 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_127_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4721__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6345_ _2338_ _2351_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6276_ _0855_ _2252_ _2287_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _1326_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4875__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6474__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _0981_ _1289_ _1291_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ _3232_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__B2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4115__I _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6162__A1 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__A1 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7238__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5976__A1 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4779__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__C _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7388__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__I _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__S _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _3372_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5900__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _0589_ _3509_ _3351_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6130_ _0960_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6456__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ _0949_ _1985_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5012_ as2650.psu\[7\] _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6208__A2 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _2941_ _2942_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5967__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ _2769_ _2873_ _2876_ _2638_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5845_ _1511_ _1437_ _1869_ _1618_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3993__A3 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5776_ _1804_ _1806_ _1807_ _1319_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4727_ _0909_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3774__I _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4942__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6144__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _0671_ _0827_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3609_ _3143_ _3144_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7377_ _0200_ clknet_leaf_12_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4589_ _0773_ _0693_ _0775_ _0715_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _1663_ _2337_ _2342_ _2266_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6447__A2 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6259_ net3 _3341_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3681__A2 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5958__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4273__C _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5186__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4933__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A1 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6135__B2 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4697__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4449__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5949__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__B2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__B1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3960_ _3288_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3891_ _3425_ _3426_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ net25 _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5561_ _1310_ _1559_ _1604_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_129_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7300_ _0123_ clknet_leaf_44_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6126__A1 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4512_ _3527_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5492_ _3233_ _1523_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7231_ _0054_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4443_ _3214_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6838__C _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7162_ _1715_ _3100_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4374_ _0395_ _0559_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4152__A3 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6113_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6429__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _3050_ _3051_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6044_ _1132_ _2059_ _2060_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4860__A1 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6946_ net39 _2925_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4612__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6877_ _3309_ _2859_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5828_ _1747_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5168__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__B2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ _1783_ _1786_ _1791_ _1759_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4915__A2 _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6117__A1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6117__B2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7429_ _0252_ clknet_leaf_3_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5425__S _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4679__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5652__C _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6840__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6108__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7426__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__A2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5134__I _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3893__A2 _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7084__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _0284_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5070__S _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6800_ _1821_ _2768_ _2785_ _1084_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ _3569_ _3504_ _0741_ _0337_ _0373_ _0490_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6731_ _3547_ _3549_ _3551_ _1533_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3943_ _3220_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6662_ as2650.addr_buff\[7\] _3235_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3874_ _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6898__A2 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _0923_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _0971_ _2584_ _2589_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ net23 _1590_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5570__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5475_ _1173_ _1524_ _1531_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6568__C _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7214_ _0037_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4426_ as2650.r123\[1\]\[7\] _0616_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5322__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7145_ _1546_ _1729_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4357_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5044__I _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3884__A2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__I1 as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7076_ _1700_ _0785_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4288_ _3563_ _0488_ _0491_ _3352_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6822__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _1989_ _2040_ _2047_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4833__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6586__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _2908_ _2905_ _2907_ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4061__A2 _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__A2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6510__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3875__A2 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6494__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3627__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6577__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_70 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_73_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_81 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_92 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6513__I _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__I as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3590_ _3125_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__A2 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5260_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4211_ _0401_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5191_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7057__A2 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ _0346_ _0290_ _0308_ _3388_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_95_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ as2650.r123\[2\]\[2\] _3451_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4815__A1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6568__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4975_ _1144_ _1102_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6714_ _1664_ _2012_ _2702_ _1672_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3926_ _3460_ _3458_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5791__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _2606_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3857_ _3392_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ as2650.stack\[7\]\[0\] _2579_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3788_ _3323_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ net22 _1574_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _1515_ _1490_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4409_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _1455_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _1132_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7048__A2 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__B1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _1009_ _3017_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7271__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__A1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5082__I1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__A1 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__B _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__A1 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5840__C _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7113__B _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6798__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5412__I _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5470__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__A2 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4028__I _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3867__I _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5773__A2 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3711_ _3246_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4691_ _3266_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _0648_ _2441_ _1030_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3642_ _3177_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6722__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5525__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6361_ _0989_ _2230_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ as2650.stack\[1\]\[7\] _1391_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6292_ _2264_ _2305_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5289__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5243_ _0706_ _1350_ _1352_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3839__A2 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__C _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5174_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4125_ _3163_ _3422_ _3564_ _3534_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6789__A1 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7294__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4056_ _3464_ _3469_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6862__B _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5213__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4016__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6153__I _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__B1 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4958_ _3507_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3775__A1 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3909_ _3400_ _3443_ _3444_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ _1052_ _1055_ _1058_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_6628_ _1907_ _2616_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ _2552_ _2564_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__B _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4255__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5452__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6491__C _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3687__I _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4007__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6063__I _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A1 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3766__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6666__C _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4246__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4981__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5930_ _1947_ _1953_ _1620_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _1885_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7069__I _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5792_ _0904_ _3227_ _3277_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6943__A1 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3757__A1 as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4743_ as2650.stack_ptr\[0\] _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4674_ as2650.psl\[7\] _0670_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6413_ _1212_ as2650.stack\[5\]\[12\] as2650.stack\[4\]\[12\] _2072_ _2426_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3625_ _3160_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7393_ _0216_ clknet_leaf_52_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6171__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4182__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _0825_ _2331_ _2358_ _2034_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4721__A3 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6275_ _2122_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7120__A1 _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__S _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5226_ _1327_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ as2650.stack\[3\]\[9\] _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4108_ _3321_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5088_ as2650.pc\[11\] _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4237__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _3563_ _3567_ _3571_ _3572_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__A2 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3748__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__I _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4131__I _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A1 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7111__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3970__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6465__A3 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__A2 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6007__B _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6925__A1 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5728__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4400__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _3508_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3911__A1 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7102__A1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6060_ _0951_ _1983_ _2081_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _0844_ _0800_ _1166_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_97_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ net39 _2674_ _1151_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5600__I _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5967__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3978__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _0936_ _0887_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7169__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6893_ _2611_ _2875_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7332__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5844_ _0922_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6916__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ _0819_ _1802_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6392__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4726_ _0316_ _0623_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4942__A3 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ _0823_ _0825_ _0831_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4155__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3608_ as2650.ins_reg\[0\] _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7376_ _0199_ clknet_leaf_12_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4588_ _0537_ _0694_ _0644_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4886__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6327_ _2264_ _2331_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3790__I _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _0939_ _1328_ _1331_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _2129_ _2207_ _2127_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6606__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4697__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3914__B _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5646__A1 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4449__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7121__B _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7355__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__A2 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__B2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4036__I _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _3409_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6251__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _1603_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_38_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ _0664_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5491_ _0760_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7230_ _0053_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4442_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _3083_ _3112_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4373_ _0402_ _0561_ _0572_ _0574_ _0395_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6200__B _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4152__A4 _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6112_ _0959_ net1 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7092_ _0453_ _3040_ _0527_ _3036_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6834__B1 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _1425_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4860__A2 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _2924_ _2902_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _2834_ _0583_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5827_ _1554_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3785__I _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1708_ _1754_ _1744_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4709_ as2650.stack_ptr\[2\] _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6117__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _1726_ _0440_ _1704_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7428_ _0251_ clknet_leaf_24_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__A2 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5876__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7359_ _0182_ clknet_leaf_27_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5240__I _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5800__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4367__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6108__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6939__C _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4842__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6044__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _1131_ _3310_ _2617_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3942_ _3402_ _3476_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ _1171_ _3486_ _3489_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_3873_ _3220_ _3249_ as2650.ins_reg\[7\] _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5612_ _3175_ _1508_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6592_ as2650.stack\[7\]\[7\] _2585_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5543_ _1149_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _1529_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5858__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7213_ _0036_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4425_ _0554_ _0615_ _0619_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7144_ _1728_ _1714_ _3097_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4356_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6865__B _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7075_ _1305_ _3014_ _3027_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4287_ _0490_ _3367_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1461_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4385__B _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5060__I _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6586__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5995__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _2908_ _2347_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_74_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6859_ _2834_ _0599_ _2842_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6338__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A1 _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5010__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A3 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__A3 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_60 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_71 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_82 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_127_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4588__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_93 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _0414_ _0295_ _0303_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4512__A1 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6685__B _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4984__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4141_ _0309_ _0310_ _3546_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ _3578_ _0278_ _3447_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6017__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6568__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6704__I _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _0914_ _3247_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_53_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3925_ as2650.holding_reg\[1\] _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6713_ _2015_ _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4224__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6644_ _2249_ _2634_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _3170_ _3172_ _3238_ _3241_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_137_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6575_ _2576_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3787_ _3167_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6740__A2 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ _0884_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ as2650.cycle\[6\] _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _3285_ _3338_ _3449_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4503__A1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5388_ as2650.stack_ptr\[1\] as2650.stack_ptr\[0\] _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7127_ _1735_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4339_ _0541_ _3367_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6256__B2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _3229_ _0802_ _1055_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_86_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6009_ _0867_ _2028_ _2031_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6008__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__B2 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7416__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A2 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6731__A2 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6798__A2 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4309__I _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5849__B _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5222__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ _3158_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3784__A2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3641_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4979__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6722__A2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5525__A3 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4733__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ _0825_ _2373_ _2034_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ _0966_ _1390_ _1394_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6291_ _1902_ _2299_ _2306_ _1572_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5289__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__A1 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5242_ as2650.r123_2\[1\]\[1\] _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5173_ _1295_ _3171_ _1296_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_96_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4124_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4055_ _3455_ _3476_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4264__A3 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4957_ _3373_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3908_ _3419_ _3399_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3775__A2 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _0829_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _1907_ _2616_ _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3839_ _3367_ _3370_ _3374_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3793__I _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _1151_ _2563_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6102__C _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5509_ _0913_ _1558_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6489_ _0751_ _0278_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6477__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4838__B _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6229__A1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6229__B2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4129__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5452__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3968__I _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A2 _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7124__B _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6640__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5443__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5860_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ as2650.pc\[10\] _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _3225_ _3226_ _3363_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3757__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4742_ _0512_ _0921_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_109_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4673_ as2650.psl\[6\] _3337_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6412_ _2415_ _2424_ _1765_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3624_ as2650.ins_reg\[2\] _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7392_ _0215_ clknet_leaf_45_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ _0855_ _2354_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6274_ _2288_ _2289_ _2290_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _1340_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5131__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5156_ _1274_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3693__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6873__B _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4107_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5087_ _1245_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6631__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ _3351_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3996__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _1431_ _1993_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4945__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3920__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5399__B as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3987__A2 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5189__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A2 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5361__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3911__A2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6249__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6310__B1 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _1167_ _1177_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6861__A1 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5416__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6613__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _2678_ _2940_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _1889_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3978__A2 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ net50 _2874_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5843_ _1107_ _0813_ _0852_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6916__A2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5774_ _1663_ _1568_ _1438_ _1805_ _1318_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7029__B _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4725_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4656_ _0833_ _0834_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3607_ _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5352__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _0541_ _0712_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7375_ _0198_ clknet_leaf_15_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ _1998_ _2340_ _0839_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6257_ as2650.addr_buff\[0\] _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6852__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ as2650.stack\[2\]\[1\] _1329_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5655__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _2171_ _2181_ _2205_ _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ as2650.stack\[3\]\[2\] _1277_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6080__A2 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4407__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4091__A1 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4918__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6778__B _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__I1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7096__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3657__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5701__I _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7020__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5582__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A2 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4510_ _3492_ _0687_ _0688_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5490_ _1541_ _1526_ _1543_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4441_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4137__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__I _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7160_ as2650.psu\[3\] _3109_ _3111_ _3096_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4372_ _0419_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7087__A1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6111_ _0960_ _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _0452_ _3040_ _3048_ _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _0338_ _2061_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6834__B2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ net38 _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4671__B _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6875_ _2835_ _2803_ _2857_ _2836_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7011__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4163__S _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5826_ _1736_ _1853_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__B1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _1788_ _1789_ _0907_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4708_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5688_ _1544_ _1718_ _0870_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ _0250_ clknet_3_2_0_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5325__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _0813_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5876__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7358_ _0181_ clknet_leaf_27_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6309_ _0855_ _2299_ _2324_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ _0112_ clknet_leaf_44_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3639__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6140__I3 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6617__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__I _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5800__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4581__B _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3811__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7002__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4367__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6301__B _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3878__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7322__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6955__C _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7132__B _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4055__A1 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4990_ as2650.psl\[7\] _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _3460_ _3475_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3802__A1 _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3886__I _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6660_ _3371_ _3390_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3872_ _3404_ _3405_ _3406_ _3407_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_108_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5611_ _1298_ _1618_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5555__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _0966_ _2584_ _2588_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _1581_ _1583_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5307__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _1522_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4424_ as2650.r123\[1\]\[6\] _0616_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7212_ _0035_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3869__A1 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4355_ as2650.holding_reg\[7\] _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7143_ _1322_ _0876_ _1729_ _0878_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4530__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6807__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6807__B2 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7074_ _1178_ _3028_ _3033_ _2736_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4286_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6025_ _2041_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A2 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _1494_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6858_ _2807_ _2810_ _2841_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5809_ _1837_ _1838_ _1575_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5546__A1 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4349__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6594__I0 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _2613_ _2774_ _1682_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5561__A4 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5849__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6775__C _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6347__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4037__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_61 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_72 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_83 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_94 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_14_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__C1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A1 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__C _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5870__B _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4512__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ _3389_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6257__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _0277_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4276__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7218__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4973_ _1143_ _3397_ _3428_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5776__B2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6712_ _1801_ _2692_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3924_ as2650.holding_reg\[1\] _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6643_ _2597_ _2607_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5528__A1 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3855_ _3390_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4200__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ _2577_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3786_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_22_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5525_ _1571_ _1573_ _0875_ _3221_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_117_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5456_ _1511_ _1512_ _1416_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4407_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4503__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5387_ _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _2249_ _3082_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4269_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _3138_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7057_ _1036_ _1019_ _3015_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6008_ _1210_ as2650.stack\[3\]\[2\] as2650.stack\[2\]\[2\] _1930_ _2030_ _2031_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6731__A3 _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__I _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6495__A2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4258__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__B1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4325__I _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6707__B1 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6707__C2 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _3173_ _3175_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6183__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6722__A3 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A4 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5156__I _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__A1 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ as2650.stack\[1\]\[6\] _1391_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6290_ _2211_ _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4995__I _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__A2 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _1348_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _0621_ _1300_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6238__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4054_ _3587_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5997__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7190__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6410__A2 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _1125_ _0871_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4421__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3907_ _3403_ _3408_ _3431_ _3442_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3775__A3 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _1054_ _1057_ _0998_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6450__I _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6626_ _1495_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6174__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3838_ _3373_ _3367_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4724__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ _0537_ _2464_ _2556_ _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3769_ _3195_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5508_ _0902_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6488_ _1154_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6477__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _0909_ _1496_ _1082_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4488__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__C _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7109_ _0823_ _0805_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5988__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5685__B _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A1 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5704__I _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__A1 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7140__B _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6640__A2 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4651__A1 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ _0981_ _0982_ _0984_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _1787_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4403__A1 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3894__I _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6156__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ _0677_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _1718_ _2423_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5903__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3623_ as2650.ins_reg\[3\] _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7391_ _0214_ clknet_leaf_45_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5903__B2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6342_ _2239_ _2355_ _2356_ _1969_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6273_ _2119_ as2650.stack\[3\]\[8\] as2650.stack\[2\]\[8\] _2241_ _2162_ _2290_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7120__A3 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ _0977_ as2650.stack\[2\]\[8\] _1327_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _1275_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3693__A2 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4106_ _3543_ _0290_ _0308_ _3300_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_99_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5086_ as2650.stack\[5\]\[10\] _1244_ _1238_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4037_ _3570_ _3563_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6631__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6445__I _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__A1 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _0943_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3748__A3 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4939_ as2650.psl\[6\] _0541_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4945__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6609_ _1420_ _1551_ _1046_ _1578_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_1_0_wb_clk_i clknet_3_4_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__B _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A3 _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6870__A2 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6622__A2 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4397__B1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__B _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6138__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7429__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7135__B _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__B2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _0989_ _2698_ _2932_ _2935_ _2936_ _2939_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4624__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _0891_ _1886_ _1890_ _1935_ _1591_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6891_ _2828_ _2832_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _1309_ _1508_ _1558_ _1420_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5773_ _1801_ _1802_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4724_ _0902_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_124_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4655_ _3261_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3606_ as2650.ins_reg\[1\] _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7374_ _0197_ clknet_leaf_11_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5352__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _3345_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6325_ _1535_ _2268_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__I _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6256_ _0869_ _2267_ _2270_ _2220_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6301__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _0892_ _1328_ _1330_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6852__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5280__S _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6187_ _1799_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3666__A2 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _0939_ _1276_ _1279_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5069_ _0964_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__I0 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6368__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5591__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5963__B _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5879__B1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7096__A2 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4606__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7251__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__A1 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4333__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4440_ _3319_ _0629_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6531__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4371_ as2650.holding_reg\[7\] _3344_ _0512_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6110_ _0953_ _0948_ _1985_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _0418_ _0422_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__A2 _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6041_ _2000_ _2002_ _2062_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ _2607_ _2922_ _2923_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4073__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6874_ _0588_ _0582_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3820__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ _1423_ _1842_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__A1 as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5022__B2 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4243__I _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5756_ _1751_ _1777_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6770__A1 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6770__B2 _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5687_ _1725_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7426_ _0249_ clknet_leaf_24_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5325__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6522__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7357_ _0180_ clknet_leaf_25_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4679__A4 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4569_ _3177_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7078__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _2122_ _2320_ _2323_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7288_ _0111_ clknet_leaf_44_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _2176_ _2254_ _2255_ _2213_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6825__A2 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3639__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__A1 _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4418__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6589__A1 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7274__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3811__A2 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6761__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6789__B _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6301__C _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3878__A2 _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6277__B1 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6808__I _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6816__A2 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4827__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5252__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3940_ _3457_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3802__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ as2650.holding_reg\[0\] _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5610_ _1309_ _1005_ _1568_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5555__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ as2650.stack\[7\]\[6\] _2585_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5541_ _1585_ _1586_ _1587_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6504__A1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7211_ _0034_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4423_ _0499_ _0615_ _0618_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3869__A2 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7142_ _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4354_ _3327_ _3334_ _3340_ _3342_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_99_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7073_ _1567_ _3031_ _3028_ _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4285_ net1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6024_ _2042_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4294__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5243__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6453__I _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6926_ _2866_ _2868_ _1492_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5794__A2 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _1164_ _0549_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5808_ _1570_ _1822_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6788_ _0871_ _0470_ _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6743__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5739_ _1573_ _1764_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ _0232_ clknet_leaf_18_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5688__B _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__B1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_62 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_73 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_84 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__B1 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__C2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6734__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5707__I _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3720__A1 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _0269_ _0275_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6670__B1 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _0914_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6973__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6711_ _1568_ _2666_ _2699_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3923_ _3457_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4007__B _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6642_ _2608_ _2630_ _2632_ _2606_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3854_ _3296_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6725__A1 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _2576_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3785_ _3320_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5617__I _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4200__A2 _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4521__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5524_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5455_ _0999_ _0924_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7150__A1 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_62_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4406_ _3285_ _3338_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5386_ as2650.stack_ptr\[1\] as2650.stack_ptr\[0\] _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _3258_ _3078_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4337_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6256__A3 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7056_ _3479_ _1026_ _1559_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4268_ _0330_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6007_ _2023_ _2029_ _1969_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4199_ _3583_ _0284_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4019__A2 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__I1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6964__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _2693_ _2890_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7312__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5519__A2 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__I _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__A3 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4258__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5455__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5207__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6955__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4430__A2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6707__B2 _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4194__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3941__A1 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7132__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _1348_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5694__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5171_ _0588_ _0678_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4122_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4053_ _3274_ _3213_ _3250_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6217__B _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5049__I1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7335__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6946__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4955_ _1109_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3906_ _3433_ _3435_ _3441_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4886_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6625_ _3267_ _3303_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3837_ _3372_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4185__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _0586_ _1854_ _2560_ _2561_ _2476_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4185__B2 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3768_ _3260_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3932__A1 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5507_ _3223_ _1556_ _1504_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6487_ _2493_ _2495_ _2496_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7123__A1 _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3699_ _3233_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _1007_ _1491_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_121_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4488__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5685__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4200__B _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5369_ _1417_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _1713_ _1696_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5437__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7039_ _2997_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6127__B _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6937__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4412__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6165__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__A1 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7114__A1 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3933__C _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7208__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7358__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5979__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4100__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__A2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__I _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4671_ _0854_ _0855_ _0809_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6156__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4071__I _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6410_ _1517_ _2417_ _2419_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3622_ _3157_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7390_ _0213_ clknet_leaf_51_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5903__A2 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3914__A1 _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6341_ _1209_ as2650.stack\[3\]\[10\] as2650.stack\[2\]\[10\] _1920_ _2356_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7105__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _2112_ as2650.stack\[1\]\[8\] as2650.stack\[0\]\[8\] _2237_ _2289_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5667__A1 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ _0972_ _1334_ _1339_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5154_ _1288_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _0309_ _0310_ _3538_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5085_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6092__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6092__B2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4036_ _3569_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4642__A2 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6919__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A2 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5987_ _0937_ _1941_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4938_ _0541_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3748__A4 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4945__A3 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__I _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6147__A2 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _3156_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6608_ _1514_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__A1 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6539_ _0772_ _2463_ _2464_ _0488_ _2478_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__A1 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4397__A1 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__B2 _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5649__A1 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7180__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4321__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7151__B _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__I _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4624__A2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5910_ _1918_ _1934_ _1800_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6890_ _2648_ _2864_ _2872_ _1855_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5841_ _1182_ _1795_ _1863_ _1866_ _1796_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5772_ _0910_ _1640_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _0903_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3605_ _3140_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7373_ _0196_ clknet_leaf_54_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4585_ _0374_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A3 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5625__I _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _2172_ _2338_ _2180_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _0975_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5206_ as2650.stack\[2\]\[0\] _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6186_ _2179_ _2194_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ as2650.stack\[3\]\[1\] _1277_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5068_ _1231_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5663__I1 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ _3393_ _3552_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6368__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A1 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5879__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6794__C _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3939__B _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__C _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _0412_ _0563_ _0571_ _0445_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _3568_ _2001_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6209__C _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6942_ net38 _2794_ _2826_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6873_ _2258_ _2854_ _2609_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6225__B _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__I _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5824_ _1423_ _1604_ _1849_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5755_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6770__A2 _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4706_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5686_ _1724_ _0396_ _1705_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7056__B _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7425_ _0248_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4637_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5355__I _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6522__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7356_ _0179_ clknet_leaf_27_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4568_ _0467_ _0709_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6895__B _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _2288_ _2321_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7287_ _0110_ clknet_leaf_44_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _0639_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6238_ _0969_ _0538_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4836__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _0489_ _2142_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3603__I _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7419__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6589__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__C _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4434__I _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__B1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6761__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5564__A3 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4772__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6277__B2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4827__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6029__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5252__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__B _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _3336_ _3292_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6201__A1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _1036_ _1307_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ as2650.addr_buff\[1\] _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5175__I _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ as2650.r123\[1\]\[5\] _0616_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7210_ _0033_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3869__A3 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7141_ _0840_ _1861_ _0843_ _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_113_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4353_ _0356_ _0554_ _0555_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6268__A1 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6268__B2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7072_ _1094_ _0423_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ _0486_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6023_ _1990_ _1992_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6925_ _2646_ _2390_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _2640_ _2838_ _2839_ _2647_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ as2650.cycle\[4\] _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6787_ _2742_ _2771_ _2743_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_3999_ _3532_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5738_ _1413_ _1765_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5669_ _1710_ _3460_ _1705_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7408_ _0231_ clknet_leaf_20_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7339_ _0162_ clknet_leaf_25_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6259__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7241__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7391__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5234__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6431__A1 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_63 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_74 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_85 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__B2 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6734__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6312__C _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6498__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__I _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3720__A2 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6670__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4276__A3 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6670__B2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__A1 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4971_ _1141_ _0580_ _1027_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6710_ _1461_ _2018_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3922_ _3356_ _3358_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6641_ _1208_ _2631_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3853_ _3386_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6725__A2 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6572_ _0895_ _0899_ _1214_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3784_ _3149_ _3319_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ _1428_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6489__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _1439_ _0913_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7150__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7264__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4405_ _0356_ _0605_ _0606_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5385_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4336_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7124_ _1723_ _3079_ _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _0671_ _1107_ _0827_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4249__I _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4267_ as2650.r0\[5\] _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6661__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5464__A2 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _2024_ as2650.stack\[1\]\[2\] as2650.stack\[0\]\[2\] _2025_ _2029_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_31_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4198_ _3426_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__I _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5216__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6413__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6413__B2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6908_ net37 _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4975__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6839_ _2819_ _2823_ _1647_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5543__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6652__A1 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5455__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A1 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6707__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4194__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6977__C _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3941__A2 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5694__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5170_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4121_ _0324_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6643__A1 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A2 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _3584_ _3585_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_84_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4954_ _0378_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3905_ _3436_ _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4885_ _0670_ _0827_ _0845_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_138_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6624_ _1487_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3836_ _3371_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4185__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5382__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3767_ _3302_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6555_ _1546_ _2522_ _1633_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5506_ _0646_ _0814_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3698_ as2650.addr_buff\[6\] _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6486_ _1856_ _3552_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6459__I _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5437_ _1492_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6331__B1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5363__I _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5685__A2 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ _0906_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7107_ _3020_ _3062_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4319_ _0512_ _0419_ _0412_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5299_ _0938_ _1384_ _1387_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__A2 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7038_ _0354_ _2998_ _3004_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__B _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4707__I _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4660__A3 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A2 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4442__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6625__A1 _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4100__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7050__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4939__A1 as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6053__B _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3611__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4670_ _0824_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3621_ _3151_ _3156_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5892__B _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3914__A2 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6340_ _2199_ as2650.stack\[1\]\[10\] as2650.stack\[0\]\[10\] _1252_ _2355_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7105__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6271_ _1457_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5222_ as2650.stack\[2\]\[7\] _1335_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5667__A2 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5153_ _0977_ as2650.stack\[3\]\[8\] _1275_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5419__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4104_ _3296_ _3360_ _3502_ _0288_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_5084_ as2650.pc\[10\] _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4890__A3 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4035_ _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A3 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6919__A2 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1616_ _1630_ _1108_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5358__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ _1035_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _0901_ _1517_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3819_ as2650.r0\[1\] _3331_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6538_ _1544_ _2522_ _1634_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _2458_ _3527_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6855__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6607__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__B _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__A1 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__A1 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5594__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A1 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5932__S _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6846__A1 _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5649__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5731__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__I1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4085__A1 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__B _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3832__A1 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _0831_ _1199_ _1865_ _1003_ _1571_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5771_ _1801_ _1658_ _1802_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__I _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _3197_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4653_ _0835_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3604_ _3139_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7372_ _0195_ clknet_leaf_40_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4584_ _0707_ _0770_ _0771_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6323_ _1989_ _2331_ _2337_ _1994_ _1753_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_89_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6837__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6837__B2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _1234_ _2221_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5205_ _1326_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _2033_ _2171_ _2198_ _2203_ _1452_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_69_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5136_ _0892_ _1276_ _1278_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5112__I1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ as2650.stack\[5\]\[5\] _1230_ _1227_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4076__A1 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__B _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ _3547_ _3549_ _3551_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_84_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5969_ _1949_ _1950_ _1991_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5088__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__A2 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6828__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4876__B _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6647__I _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4167__I _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5103__I1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4067__A1 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5803__A2 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5726__I _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6819__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6295__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6047__A2 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4058__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6941_ _1244_ _2637_ _2921_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _2258_ _2854_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_90_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ _1850_ _0833_ _1719_ _1818_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_124_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5754_ _1516_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_56_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4230__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_120_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5685_ _1541_ _1697_ _1723_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7424_ _0247_ clknet_leaf_31_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4636_ _3178_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7355_ _0178_ clknet_3_3_0_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4533__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5730__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _0686_ _0754_ _0755_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6895__C _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6306_ as2650.stack\[7\]\[9\] _1455_ _2241_ as2650.stack\[6\]\[9\] _2074_ _2322_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7286_ _0109_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4498_ _0634_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6467__I _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6237_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5371__I _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6168_ _1894_ _2182_ _2186_ _1718_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5119_ as2650.stack\[4\]\[8\] _1237_ _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _2119_ as2650.stack\[3\]\[4\] as2650.stack\[2\]\[4\] _1929_ _1468_ _2120_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_100_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5797__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4715__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6135__C _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5549__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6746__B1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__B2 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A1 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4072__I1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5564__A4 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5990__B _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4827__A3 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5788__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__B _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4460__A1 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__C _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6201__A2 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7157__B _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5470_ _1487_ _1524_ _1527_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4421_ _0424_ _0615_ _0617_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7140_ _1165_ _0877_ _1810_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4352_ as2650.r123\[2\]\[6\] _0425_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4283_ _3164_ _0359_ _0457_ _0448_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ _2539_ _2540_ _3030_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6022_ _2043_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7193__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _2858_ _2860_ _1747_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _1136_ _2640_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5806_ _1795_ _3277_ _1832_ _1836_ _1796_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6786_ _0376_ _0388_ _0390_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4203__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3998_ _3497_ _3500_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5737_ _1426_ _1767_ _1769_ _1670_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__5951__B2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _1173_ _1643_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ _0230_ clknet_leaf_36_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4619_ _0803_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5599_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _0161_ clknet_leaf_34_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6259__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ _0092_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6431__A2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_75 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_86 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4993__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6195__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6734__A3 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5942__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_1_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5879__C _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4681__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6056__B _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6422__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _0567_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _3399_ _3455_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _1145_ _1645_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3852_ as2650.addr_buff\[5\] _3387_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__6725__A3 _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5933__A1 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A2 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _1150_ _2565_ _2575_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4304__B _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3783_ _3177_ _3318_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5522_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6489__A2 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5453_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4404_ as2650.r123\[2\]\[7\] _0425_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5384_ _1439_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7123_ _3073_ _3074_ _3075_ _3076_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4335_ net2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7054_ _1566_ _0854_ _1653_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4266_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ as2650.stack\[6\]\[2\] _1930_ _1922_ _2022_ _2027_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6661__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _3403_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ net50 _2874_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _1232_ _2665_ _2822_ _2623_ _1582_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6177__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__B2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__I0 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4727__A2 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _2658_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__A3 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6168__B2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6323__C _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4718__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5734__I _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6340__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6340__B2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__A2 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ _3336_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6643__A2 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4051_ _3459_ _3463_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 io_in[5] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A1 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4953_ _1096_ _1117_ _1122_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6514__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4813__I _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3904_ _3274_ _3439_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4884_ _1054_ _1011_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6623_ _3391_ _2613_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7231__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3835_ net5 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5906__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5906__B2 _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _2516_ _1141_ _2559_ _1138_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3766_ _3296_ _3301_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _1033_ _1045_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6485_ _2494_ _3545_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3697_ as2650.addr_buff\[5\] _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7381__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7123__A3 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _3305_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__B2 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6882__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5367_ _1424_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7106_ _1755_ _3063_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4318_ _0261_ _0516_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5298_ as2650.stack\[1\]\[1\] _1385_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6095__B1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ as2650.r123\[0\]\[3\] _3000_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6634__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4249_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__B1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6398__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6143__C _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6625__A2 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7254__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4939__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4633__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3611__A2 _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _3152_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6270_ as2650.stack\[6\]\[8\] _2195_ _1922_ _2284_ _2286_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6313__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _0967_ _1334_ _1338_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6864__A2 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _0972_ _1282_ _1287_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6509__B _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _3369_ _3564_ _3534_ _3561_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_110_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__I _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3712__I as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _1242_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ net7 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7041__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5985_ _1427_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4936_ _0757_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _1036_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6606_ net28 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ as2650.r123\[1\]\[1\] as2650.r123_2\[1\]\[1\] _3288_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6552__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ as2650.pc\[8\] _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7075__B _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6537_ _1159_ _2541_ _2543_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3749_ _3284_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3756__I3 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6468_ _1082_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6855__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ as2650.r123_2\[0\]\[3\] _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6399_ _1247_ _1243_ _2344_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4866__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6607__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3622__I _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4618__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7277__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4094__A2 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7032__A2 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5594__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7099__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4609__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__B1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5887__C _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3832__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7023__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _0904_ _3227_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4721_ _3225_ _0904_ _3224_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6534__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3603_ _3138_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7371_ _0194_ clknet_leaf_38_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ as2650.r123_2\[2\]\[5\] _0738_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3899__A2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6322_ _2333_ _2336_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4560__A3 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6298__B1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6837__A2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6253_ _1915_ _2269_ _1441_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4848__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5204_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6184_ _2159_ _2202_ _2122_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ as2650.stack\[3\]\[0\] _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4982__B _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__A1 _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ _3550_ _3535_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3823__A2 _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7014__A2 _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__I _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5968_ as2650.pc\[1\] _3505_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6773__A1 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4206__C _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4919_ _0452_ _0527_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5899_ _0898_ as2650.stack\[5\]\[0\] as2650.stack\[4\]\[0\] _0929_ _1924_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3818__S _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6525__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6421__C _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4839__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4067__A2 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5803__A3 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3814__A2 _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7005__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6819__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3750__A1 _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6059__B _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4358__I as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__A2 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6573__I _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6940_ _2916_ _2920_ _1647_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _2254_ _2817_ _2213_ _2255_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__B2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ _1572_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5753_ _1094_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6522__B _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4821__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _0363_ _1719_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7423_ _0246_ clknet_leaf_4_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4635_ _0805_ _0816_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _0177_ clknet_leaf_27_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ as2650.r123_2\[2\]\[4\] _0738_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4977__B _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5730__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6305_ _2112_ as2650.stack\[5\]\[9\] as2650.stack\[4\]\[9\] _2237_ _2321_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6748__I _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7285_ _0108_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _0319_ _0638_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6236_ _2173_ _2212_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4297__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4268__I _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6167_ _1187_ _1812_ _1007_ _3387_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5118_ _1255_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6098_ _0893_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__B _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6483__I _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5049_ as2650.stack\[5\]\[0\] _1208_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__A1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6746__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__A2 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__B2 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5827__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6432__B _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7171__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__I _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__A1 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5562__I _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4288__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4532__I0 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6594__S _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5788__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6985__A1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6342__B _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4212__A2 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__I _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7162__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ as2650.r123\[1\]\[4\] _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4351_ _3453_ _0528_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5472__I _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7070_ _0804_ _3029_ _1726_ _0808_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4282_ _0483_ _0372_ _0484_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4279__A2 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _0941_ net7 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6425__B1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4816__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7338__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6976__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6976__B2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _2612_ _2903_ _1847_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _2834_ _0582_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net13 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5805_ _1833_ _1835_ _1737_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6785_ _0388_ _0390_ _0375_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3997_ _3287_ _3530_ _3531_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5400__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _1295_ _1508_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7153__A1 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5667_ _3493_ _1708_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7406_ _0229_ clknet_leaf_37_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4618_ _0798_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5598_ _1296_ _3279_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6900__A1 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7337_ _0160_ clknet_leaf_30_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4549_ as2650.r123_2\[2\]\[3\] _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7268_ _0091_ clknet_leaf_46_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6219_ _1251_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7199_ _0022_ clknet_leaf_6_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_54 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_65 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A2 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7424__D _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__I _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7012__I _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6958__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ _3269_ _3360_ _3454_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3851_ as2650.addr_buff\[6\] _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5467__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _2568_ _2570_ _2574_ _2476_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_73_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3782_ _3251_ _3256_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5933__A2 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A3 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ _1036_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7135__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6800__B _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _1414_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4403_ _3453_ _0577_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5383_ _1411_ _1450_ _1451_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7122_ _3072_ _0875_ _0805_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4334_ _0484_ _0487_ _0529_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5449__A1 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7053_ _1541_ _3011_ _3013_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4265_ _0346_ _0372_ _0460_ _0389_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4121__A1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _2023_ _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6661__A3 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4196_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6949__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _2648_ _2886_ _2887_ _1827_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _2666_ _2178_ _2821_ _2626_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6177__A2 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6768_ _2746_ _2747_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3935__A1 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5719_ _1461_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7126__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6699_ _1534_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4230__B _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4360__A1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5045__C _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4112__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__A2 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3926__A1 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7117__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7183__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A1 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4103__A1 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4050_ _3583_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5851__A1 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[6] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5603__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _3223_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3903_ _3421_ _3438_ _3411_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4883_ _0646_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6622_ _1420_ _3236_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3834_ _3162_ _3369_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3917__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _1098_ _0448_ _2558_ _1096_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7108__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3765_ _3298_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5504_ _1017_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4590__A1 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6484_ _1682_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3696_ _3211_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5435_ as2650.cycle\[6\] _3196_ _1489_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6331__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _1423_ _1430_ _1434_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4317_ _0261_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7105_ _3193_ _1715_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5297_ _0891_ _1384_ _1386_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ _0279_ _2998_ _3003_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _0395_ _0431_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5842__B2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4179_ _3353_ _0374_ _0383_ _3323_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__S _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4948__A3 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3908__A1 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__A2 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4581__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4884__A2 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6561__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6313__A2 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4324__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ as2650.stack\[2\]\[6\] _1335_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5151_ as2650.stack\[3\]\[7\] _1283_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6077__A1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4102_ _3540_ _0288_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_116_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ as2650.stack\[5\]\[9\] _1241_ _1238_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5824__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4033_ _3503_ _3566_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6525__B _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _2004_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _1099_ _1102_ _1104_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _0757_ _1028_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6605_ _0994_ _2591_ _2596_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3817_ _3352_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4797_ _0972_ _0956_ _0973_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6552__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__A1 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3748_ _3169_ _3244_ _3257_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6536_ as2650.psl\[5\] _0848_ _2542_ _0808_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3679_ _3209_ _3212_ _3213_ _3214_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6467_ _2454_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ _1474_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6398_ _2403_ _2401_ _2410_ _1452_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4866__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5349_ _0817_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5390__I _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4079__B1 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4618__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _2961_ _0785_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5291__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4734__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4554__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__I _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6059__A1 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4609__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__B2 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7371__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5585__A3 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4720_ as2650.cycle\[2\] _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _3224_ _3154_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6534__A2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3602_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4545__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7370_ _0193_ clknet_leaf_39_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4582_ _0453_ _0752_ _0756_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_122_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6321_ _2334_ _2335_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6252_ _1525_ _2268_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6298__B2 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4848__A2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6183_ _2110_ _2200_ _2201_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3723__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5134_ _1274_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ as2650.pc\[5\] _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4982__C _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _3546_ _3548_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6470__A1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6222__B2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ as2650.pc\[2\] net7 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4784__A1 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4918_ _0422_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5898_ as2650.stack\[7\]\[0\] _1465_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_139_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ _0409_ _1017_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6525__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5385__I _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _2494_ _0362_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6289__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4839__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6944__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7394__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5264__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6461__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__I _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5972__B1 _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5295__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3808__I _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__A2 _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4527__A1 _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3750__A2 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4639__I _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5255__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6870_ _2828_ _2678_ _2853_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5007__A2 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ _1845_ _1846_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6755__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4215__B1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5752_ _1453_ _1780_ _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4703_ as2650.pc\[0\] _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _1722_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3718__I _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7422_ _0245_ clknet_leaf_6_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4042__C _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7267__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7353_ _0176_ clknet_leaf_35_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4565_ _0749_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6304_ _2239_ _2318_ _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7284_ _0107_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4496_ _0662_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6235_ _0974_ _2251_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_103_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6691__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6166_ _1052_ _2183_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _1265_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6097_ _2024_ as2650.stack\[1\]\[4\] as2650.stack\[0\]\[4\] _2025_ _2118_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5048_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _2969_ _2974_ _2975_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6746__A2 _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__A1 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3628__I _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3980__A2 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3732__A2 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4459__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6682__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6682__B2 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__B _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4996__A1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4922__I _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6342__C _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7162__A2 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4350_ _3485_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4920__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _3164_ _0359_ _0457_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4279__A3 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6020_ _0947_ _0337_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__I _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5228__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A2 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ net38 _2902_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6853_ _2835_ _2803_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6728__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5804_ _1421_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6784_ _0872_ _2684_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ as2650.r123\[2\]\[1\] _3451_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5735_ _1295_ _0839_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3962__A2 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ _1707_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7153__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ _0228_ clknet_leaf_37_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5164__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4617_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5597_ _1638_ _1641_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6900__A2 _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _0159_ clknet_leaf_27_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4911__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4548_ _0683_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _0090_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4479_ _3337_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6218_ _1869_ _2229_ _2235_ _2008_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7198_ _0021_ clknet_leaf_5_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6149_ _2129_ _2168_ _2127_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6416__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6416__B2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_55 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_88 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7432__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3953__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7144__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5573__I _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5458__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__A1 _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__A1 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ _3385_ as2650.addr_buff\[6\] _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3781_ _3316_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5520_ _1550_ _1565_ _1569_ _1473_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7135__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6800__C _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _0835_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5483__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4601__B _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6894__A1 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4402_ _3485_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5697__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5382_ _1411_ _1450_ _0885_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7121_ _3072_ _1697_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4333_ as2650.r0\[6\] _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6646__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4264_ _3548_ _0461_ _0464_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7052_ _1567_ _3011_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__A3 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _2024_ as2650.stack\[5\]\[2\] as2650.stack\[4\]\[2\] _2025_ _2026_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4121__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4195_ _0398_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3731__I _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6949__A2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7071__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5621__A2 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _1529_ _2869_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4562__I _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6836_ _1126_ _2139_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4188__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _2682_ _2752_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3979_ _3510_ _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5718_ _1741_ _1744_ _1745_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__3935__A2 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6698_ _2652_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _3234_ _1690_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3699__A1 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4230__C _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7319_ _0142_ clknet_leaf_53_wb_clk_i as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6637__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4737__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__I _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4179__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5376__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3926__A2 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7117__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3816__I _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7328__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4351__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6628__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6348__B _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4647__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[7] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7053__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6800__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4951_ _0587_ _1120_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4382__I as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3902_ _3437_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4882_ _0641_ _3165_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ _2611_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3833_ _3368_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3917__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6552_ _0997_ _2469_ _2557_ _1652_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7108__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3764_ _3203_ _3299_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _0837_ _1551_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3726__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _1436_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3695_ _3172_ _3223_ _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6867__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5434_ _3239_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5365_ _1412_ _1432_ _1433_ _0917_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_99_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6619__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4985__C _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7104_ _0637_ _1555_ _3022_ _3025_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_141_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4316_ _0501_ _3271_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ as2650.stack\[1\]\[0\] _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6095__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7035_ as2650.r123\[0\]\[2\] _3000_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4247_ _3403_ _0432_ _0446_ _0450_ _3400_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4178_ _0378_ _3509_ _3376_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__A4 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6819_ _1164_ _0535_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3908__A2 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6858__A1 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__A2 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5800__B _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5349__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6849__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4324__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5761__I _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _0967_ _1282_ _1286_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6078__B _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6077__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4088__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5824__A2 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4032_ _3369_ _3564_ _3511_ _3565_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_96_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5588__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _2005_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4934_ _0636_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5001__I _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4865_ as2650.halted _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6604_ as2650.stack\[7\]\[12\] _2592_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _3351_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4796_ as2650.stack\[6\]\[7\] _0957_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ as2650.psu\[5\] _2467_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5760__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3747_ _3258_ _3282_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4563__A2 _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _1650_ _2456_ _2477_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3678_ _3157_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5417_ _0723_ _1477_ _1480_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4315__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__I _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ _1899_ _2409_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _0676_ _1297_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4079__A1 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ _0971_ _1369_ _1374_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4079__B2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _2983_ _2989_ _2990_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7017__A1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5112__S _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6435__C _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6240__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6528__B1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4750__I _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4003__A1 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5751__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6677__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__A3 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__I _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5806__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4925__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5019__B1 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6231__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3985__B _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5990__A1 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4650_ _3174_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 wb_rst_i net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3601_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5742__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _0766_ _0768_ _0752_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _2259_ _2302_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6251_ _3281_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5491__I _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5202_ _0930_ _1273_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ as2650.stack\[7\]\[6\] _2115_ _1971_ as2650.stack\[6\]\[6\] _2201_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5064_ _1228_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _3548_ _3540_ _3541_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__7196__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6470__A2 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4481__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6222__A2 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5966_ _1901_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4917_ _0307_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4784__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _1466_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5666__I _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _3159_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4779_ _0955_ _0956_ _0958_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6518_ _0363_ _2509_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5615__B _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _1760_ _3446_ _2457_ _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__S _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4745__I _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6461__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4472__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5567__A4 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5972__B2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5724__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3824__I _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__B _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5820_ _3202_ _3241_ _1847_ _1603_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4215__A1 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5751_ _1642_ _0863_ _1762_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5486__I _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4702_ _0865_ _0882_ _0886_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5682_ _1721_ _0287_ _1705_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7421_ _0244_ clknet_leaf_6_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7352_ _0175_ clknet_leaf_34_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _0423_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3821__S0 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _2119_ as2650.stack\[3\]\[9\] as2650.stack\[2\]\[9\] _2241_ _1468_ _2319_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7283_ _0106_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7353__D _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3734__I _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _0631_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6234_ _0970_ _2209_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6691__A2 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _1431_ _2171_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ as2650.stack\[4\]\[7\] _1235_ _1261_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6266__B _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _1469_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5047_ _0899_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_34_wb_clk_i clknet_opt_2_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4454__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4206__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6998_ net42 _2970_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7097__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5949_ _0897_ as2650.stack\[1\]\[1\] as2650.stack\[0\]\[1\] _1972_ _1973_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7211__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7361__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__A2 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5173__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4920__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _3183_ _3275_ _0357_ _0462_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A2 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6921_ net37 net50 _2874_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _1164_ _0534_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6728__A3 _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _1135_ _1000_ _1500_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7234__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _1606_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5936__A1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ _3453_ _3484_ _3529_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _0921_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _1105_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7384__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _0227_ clknet_leaf_37_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4616_ _3436_ _0645_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6361__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7335_ _0158_ clknet_leaf_24_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4911__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ _0307_ _0627_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7266_ _0089_ clknet_leaf_48_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4478_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6217_ _1137_ _2059_ _2005_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7197_ _0020_ clknet_leaf_5_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5872__B1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _2131_ _2138_ _2167_ _2037_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _1894_ _2095_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4427__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_56 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_14_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6352__A1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__B2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6655__A2 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6407__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7257__CLK clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7080__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A2 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3780_ as2650.r0\[0\] _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6591__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5764__I _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5450_ _3278_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5146__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _3315_ _0583_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6894__A2 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5381_ _1449_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7120_ _3073_ _3074_ _3075_ _3076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4332_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6809__B _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6646__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__A3 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7051_ _1537_ _3011_ _3012_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4263_ _0455_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4657__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _1211_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5854__B1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6528__C _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4194_ _0396_ _0397_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_67_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5004__I _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7071__A2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _1529_ _2861_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6835_ _2667_ _2797_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5909__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ _0378_ _3267_ _2647_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3978_ _3164_ _3437_ _3512_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5717_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6697_ _3570_ _3552_ _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6334__A1 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5648_ _1689_ _1691_ _1692_ _1473_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5137__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5932__I1 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5579_ _3210_ _3188_ _3370_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__3699__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4896__A1 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7318_ _0141_ clknet_leaf_53_wb_clk_i as2650.stack_ptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6637__A2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _0072_ clknet_leaf_46_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7062__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__B1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4753__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5376__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6325__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6876__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5533__B _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4928__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 io_in[8] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3862__A2 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__I _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6800__A2 _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _1095_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3901_ _3416_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4881_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5695__S _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6013__B1 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6620_ _1493_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3832_ _3291_ _3293_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6564__A1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ net27 _0847_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3763_ as2650.idx_ctrl\[0\] _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5494__I _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5502_ _3397_ _3221_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6316__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _1713_ _2455_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3694_ _3209_ _3229_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5433_ _0906_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6867__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _1051_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7422__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7103_ _1582_ _0559_ _3060_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6619__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4315_ _3271_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _1382_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _3530_ _2998_ _3002_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4246_ _0447_ _0449_ _0301_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ _3508_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3853__A2 _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A2 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__B _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _2777_ _2801_ _2802_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6555__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6749_ _2707_ _2678_ _2735_ _2736_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6307__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__A2 _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6449__B _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__I _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3652__I as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5669__I0 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4097__A2 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7035__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5046__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6184__B _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A2 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6912__B _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6546__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5349__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6849__A2 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ _0281_ _0284_ _0302_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_123_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ as2650.pc\[9\] _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4088__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5285__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ _3163_ _3369_ _3564_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6806__C _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7026__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5037__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6785__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5588__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _3156_ _0924_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3599__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _1103_ _1099_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4864_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6537__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _0990_ _2591_ _2595_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3815_ _3149_ _3350_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3737__I _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4795_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4012__A2 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_59_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6534_ _2539_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _3265_ _3276_ _3281_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_107_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6465_ _2461_ _2475_ _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3677_ _3188_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5416_ as2650.r123_2\[0\]\[2\] _1478_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6396_ _2407_ _2408_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5347_ _1414_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5278_ as2650.stack\[0\]\[7\] _1370_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7017_ net19 _2986_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4229_ _0429_ _0430_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7318__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6776__A1 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4251__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6528__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__B2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3647__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A1 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4003__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__B2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5751__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__A1 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__I _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6693__I _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7008__A2 _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__A1 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4490__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__B2 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4146__C _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__C _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5990__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3600_ as2650.psl\[4\] _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4580_ _0470_ _0767_ _0703_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5742__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6250_ _1432_ _2252_ _2265_ _2266_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6298__A3 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _1325_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6181_ _2111_ as2650.stack\[5\]\[6\] as2650.stack\[4\]\[6\] _2199_ _2200_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5132_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5258__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ as2650.stack\[5\]\[4\] _1226_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6536__C _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4014_ _3488_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6758__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5965_ _1896_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4233__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4851__I _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4916_ _3446_ _1086_ _0278_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5896_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4847_ _3219_ _0646_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6930__A1 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ as2650.stack\[6\]\[4\] _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6930__B2 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3744__A1 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3729_ _3260_ _3264_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6517_ _1650_ _2508_ _2525_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _1827_ _3391_ _2459_ _1768_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4298__I as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6379_ _1426_ _2373_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__S _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4472__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7290__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4761__I _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5972__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7174__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6516__A4 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6921__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6688__I _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__I _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4936__I _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3840__I _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6988__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A2 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4215__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5750_ _1777_ _1778_ _1781_ _1782_ _1453_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ as2650.psu\[5\] _0865_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5681_ _1537_ _1697_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7165__B2 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7420_ _0243_ clknet_leaf_8_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4632_ _0678_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5715__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6912__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7351_ _0174_ clknet_3_4_0_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4563_ _3258_ _3265_ _3276_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_116_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3821__S1 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _2112_ as2650.stack\[1\]\[9\] as2650.stack\[0\]\[9\] _2237_ _2318_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7282_ _0105_ clknet_leaf_3_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4494_ _0684_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6233_ _1798_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1662_ _2178_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5115_ _1264_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6039__S _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ as2650.stack\[7\]\[4\] _2115_ _1971_ as2650.stack\[6\]\[4\] _2116_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6979__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6266__C _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1210_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__B _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4454__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6997_ _2960_ _1118_ _2973_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4206__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _0927_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7156__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5879_ _1898_ _1900_ _1903_ _0889_ _1462_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6903__A1 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4390__A1 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4142__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__B2 _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5361__B _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4756__I _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__B1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6434__A3 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5642__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5587__I _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3708__A1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3835__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__A3 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7186__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4133__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5633__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6920_ _2900_ _2901_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _0540_ _0534_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5497__I _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _1512_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _2133_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3994_ _3485_ _3522_ _3528_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5936__A2 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7138__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6830__B _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ _1706_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7403_ _0226_ clknet_leaf_37_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4615_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5595_ _1609_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6361__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7334_ _0157_ clknet_leaf_17_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4546_ _0626_ _0734_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4477_ _3332_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7265_ _0088_ clknet_leaf_57_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6216_ _1812_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7196_ _0019_ clknet_leaf_5_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__B2 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _2137_ _2158_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _2096_ _2098_ _2018_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _0584_ _1105_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_57 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_79 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3938__A1 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7127__I _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__I _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6915__B _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A1 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6591__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _3313_ _0597_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5380_ _1413_ _1422_ _1435_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ _0454_ _0530_ _0531_ _0456_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4597__S _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5780__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4106__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7050_ _1573_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4106__B2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4262_ _0456_ _0460_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6001_ _1251_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4657__A2 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5854__B2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ _0396_ _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6949__A4 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6544__C _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ _2607_ _2884_ _2885_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5621__A4 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _2798_ _2815_ _2818_ _1857_ _2457_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7351__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5909__A2 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6765_ _2748_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6582__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3977_ _3296_ _3511_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5716_ _1748_ _1749_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4593__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6696_ _1172_ _3490_ _3491_ _2650_ _2651_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_136_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ _3299_ _1689_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__B2 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _0874_ _0829_ _1622_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_89_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4896__A2 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7317_ _0140_ clknet_leaf_53_wb_clk_i as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4529_ _3552_ _0719_ _0662_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7248_ _0071_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7179_ _0002_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4255__B _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6026__I _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4584__A1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4103__A4 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 io_in[9] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_92_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7374__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3900_ _3191_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4880_ _0999_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3831_ _3366_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6564__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4575__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3762_ _3297_ _3204_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6550_ _1741_ _0528_ _2479_ _2555_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5501_ _1510_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3693_ _3224_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6481_ _3494_ _2476_ _2491_ _1695_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5432_ _3195_ _1488_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5363_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__C _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _1085_ _3038_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _0474_ _0475_ _0477_ _0479_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5294_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7033_ as2650.r123\[0\]\[1\] _3000_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4245_ _0440_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5015__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4176_ _0329_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6555__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__I _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6004__A1 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6817_ _2799_ _2800_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4566__A1 as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ _1472_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ _1129_ _2667_ _2668_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4318__A1 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7247__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5669__I1 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6491__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5809__B _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5595__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5544__B _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5036__S _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ _3458_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5285__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6482__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5824__A4 _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5981_ _2000_ _2002_ _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6785__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5588__A3 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3599__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ _0536_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ as2650.stack\[7\]\[11\] _2592_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3814_ _3192_ _3349_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4794_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _2465_ _0482_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3745_ _3280_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4563__A4 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _2454_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3676_ _3211_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ _0706_ _1477_ _1479_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6395_ as2650.pc\[12\] _0540_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5346_ _3197_ _0905_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5277_ _0966_ _1369_ _1373_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6473__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7016_ _0471_ _2976_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4228_ _0430_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ _0320_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6225__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5028__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A3 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5200__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4759__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6700__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A3 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4494__I _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6216__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6923__B _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6642__C _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5200_ _1026_ _1303_ _1311_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _1211_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _1214_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5062_ _1216_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4013_ _3536_ _3537_ _3546_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6758__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _1985_ _1986_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6552__C _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ _3456_ _3482_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4846_ _3232_ _3177_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _0931_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3744__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4941__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6516_ _2509_ _2514_ _2515_ _2524_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_3728_ _3263_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__I _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6447_ _2458_ _3303_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3659_ as2650.cycle\[7\] _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6694__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _2389_ _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5329_ _1404_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5249__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6997__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5203__I _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4247__C _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7435__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6749__A2 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__B _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3680__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__C _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3658__I _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3983__A2 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5806__C _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6685__A1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6918__B _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5314__S _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6437__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4952__I _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4700_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _0725_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5176__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6373__B1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7350_ _0173_ clknet_leaf_11_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4562_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _1655_ _2314_ _2316_ _1940_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_143_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7281_ _0104_ clknet_leaf_3_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4493_ _0685_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6220__S0 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6232_ _1735_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6163_ _0965_ _2148_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5224__S _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5114_ as2650.stack\[4\]\[6\] _1232_ _1261_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _1455_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6979__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6119__I _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _0920_ _0926_ _1213_ _3264_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4067__C _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _3494_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5403__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5947_ _1919_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5167__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4390__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7479_ net46 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__B _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6419__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__C _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A1 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7092__B2 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__A2 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7147__A2 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5158__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4905__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5173__A4 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5552__B _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4133__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4947__I _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5881__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7083__A1 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4841__B1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5778__I _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4682__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6850_ net3 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _1637_ _1830_ _1831_ _1567_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6781_ _2134_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3993_ _3245_ _3311_ _3527_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5732_ _3246_ _1616_ _1629_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7138__A2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5663_ _1699_ _3407_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7402_ _0225_ clknet_leaf_37_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6897__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4614_ _3180_ _3182_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ _1043_ _1640_ net53 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7333_ _0156_ clknet_leaf_17_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4545_ _0313_ _0703_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6649__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7264_ _0087_ clknet_leaf_57_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4476_ _3446_ _0627_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7280__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6215_ _1135_ _3341_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5321__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _0018_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6146_ _1429_ _2131_ _2165_ _1927_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6077_ _2053_ _2083_ _2097_ _1810_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6821__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5624__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5028_ _1161_ _1156_ _0804_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_input10_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_58 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ net40 _2674_ _0885_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4060__A1 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6888__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4363__A2 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4767__I _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__A1 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3671__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7065__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6812__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5615__A2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3626__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5551__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4330_ _3523_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4106__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5303__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _3523_ _0461_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _1974_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5854__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ _0324_ _0326_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3865__A1 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7056__A1 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6803__A1 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ net50 _2794_ _2826_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6833_ _2173_ _2817_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6764_ _2749_ _2750_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ as2650.ins_reg\[4\] _3275_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4042__A1 _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5715_ _1548_ _1636_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4593__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _2653_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5646_ _3233_ _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5542__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5577_ _0876_ _3319_ _1037_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5971__I _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7316_ _0139_ clknet_leaf_64_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ _0631_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7247_ _0070_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4459_ _0650_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7178_ _0001_ clknet_leaf_3_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3856__A1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _1225_ _2094_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4281__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4033__A1 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4887__A3 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5836__A2 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__B _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7038__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6261__A2 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4272__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__C _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A2 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4960__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3830_ _3148_ _3365_ _3222_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4024__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3761_ as2650.idx_ctrl\[1\] _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5772__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ net24 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _2478_ _2483_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3692_ _3225_ _3226_ _3227_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_118_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _3154_ _3279_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4878__A3 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5362_ _0677_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _3346_ _3034_ _3059_ _2736_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4313_ _0505_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__I1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5293_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7032_ _3448_ _2998_ _3001_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4244_ _0428_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3838__A1 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7029__A1 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7199__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4175_ _0331_ _0289_ _0379_ _3511_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5966__I _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _2799_ _2800_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4015__A1 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _2705_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6960__B1 _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3959_ _3493_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6678_ _1768_ _2639_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5515__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _0900_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4110__I as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3829__A1 _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6491__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4780__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5054__I0 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5506__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6500__I _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7341__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4020__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4955__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5052__S _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _2000_ _2002_ _0750_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4245__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _1100_ _1101_ _0584_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4796__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5993__A1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4690__I _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4862_ _0835_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ _0986_ _2591_ _2594_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3813_ _3207_ _3176_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5745__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _2471_ _0586_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3744_ _3278_ _3279_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _2462_ _2463_ _2464_ _3370_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3675_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ as2650.r123_2\[0\]\[1\] _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _2335_ _2404_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0903_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ as2650.stack\[0\]\[6\] _1370_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6566__B _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7015_ _2961_ _0772_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4865__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ _0429_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6473__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ as2650.r0\[4\] _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4086__B _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _3459_ _3463_ _0272_ _0273_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5984__A1 _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7214__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3944__I _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7364__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6476__B _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4775__I _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5975__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _1272_ _1253_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4466__A1 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4012_ as2650.addr_buff\[5\] _3387_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7237__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5963_ _0937_ _0889_ _0943_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _0576_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5894_ _1456_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5718__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _3266_ _3319_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7387__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4776_ _0932_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6930__A3 _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6515_ _0365_ _1854_ _2521_ _2523_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3727_ _3261_ _3262_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6446_ _1682_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6143__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3658_ _3185_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6143__B2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ _2279_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3589_ as2650.ins_reg\[1\] _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5328_ as2650.r123\[3\]\[1\] _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5259_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4457__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4209__A1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__C _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3680__A2 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5709__A1 _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6382__A1 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6382__B2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7146__I _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3674__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6050__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6685__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4696__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6437__A2 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4448__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _0673_ _0802_ _0809_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_124_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5176__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6373__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__B2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _0624_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _2060_ _2315_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7280_ _0103_ clknet_leaf_66_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4492_ _0669_ as2650.r123_2\[2\]\[0\] _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6231_ _0972_ _1936_ _2248_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6220__S1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6828__C _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _2172_ _2179_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__A2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5113_ _1263_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _2110_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5304__I _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5939__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6995_ _2959_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ as2650.stack\[7\]\[1\] as2650.stack\[4\]\[1\] as2650.stack\[5\]\[1\] as2650.stack\[6\]\[1\]
+ _0928_ _0897_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4611__A1 as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _0836_ _3227_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5167__A2 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ as2650.pc\[2\] _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _0679_ _1010_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__C _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4850__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6355__A1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4905__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__A1 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6929__B _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3892__A2 as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6664__B _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4963__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__B2 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5800_ _0909_ _0919_ _1824_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6780_ _2086_ _2737_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ _3525_ _3526_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5731_ _1300_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7138__A3 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6346__A1 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5149__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6346__B2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7401_ _0224_ clknet_leaf_36_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4613_ _3333_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6897__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _0155_ clknet_3_3_0_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4544_ _0349_ _0687_ _0688_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6839__B _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__CLK clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__A2 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7263_ _0086_ clknet_leaf_51_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _0666_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _2189_ _2190_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7194_ _0017_ clknet_leaf_1_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5321__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _2159_ _2160_ _2164_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5872__A3 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5034__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7074__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6076_ _1431_ _2091_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6821__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _0803_ _1195_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6293__C _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4832__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_59 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6034__B1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__A2 as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ _1690_ _2952_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _1948_ _1938_ _1952_ _1051_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4060__A2 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6337__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6337__B2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3952__I _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7065__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4783__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3626__A2 as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5379__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5551__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__I _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4191_ as2650.holding_reg\[4\] _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7056__A2 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4693__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6803__A2 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6901_ _0976_ _2636_ _2878_ _2608_ _2883_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4290__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6832_ _2175_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6763_ _2712_ _0312_ _2679_ _2713_ _2714_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3975_ _3475_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5090__I1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ _3202_ _3251_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6694_ _1130_ _2682_ _2648_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5645_ _1646_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _1585_ _1587_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7315_ _0138_ clknet_leaf_62_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4527_ _3554_ _0710_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7246_ _0069_ clknet_leaf_57_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4458_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4089__B _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ _0000_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5845__A3 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4389_ _3343_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7047__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6128_ _1229_ _1224_ _2094_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6059_ _1984_ _2080_ _1575_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4281__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5230__A1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5781__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5533__A2 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6730__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3682__I as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7038__A2 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4219__S _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6797__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__A1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7270__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3857__I _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5221__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5772__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3783__A1 _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3691_ _3152_ _3150_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_125_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _3196_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4688__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _1425_ _1426_ _1427_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3592__I _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4878__A4 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _0400_ _0407_ _0433_ _0514_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7100_ _3053_ _3054_ _3058_ _1759_ _3034_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_82_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5292_ _1214_ _1360_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ as2650.r123\[0\]\[0\] _3000_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4243_ _3274_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7029__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4174_ _3540_ _0289_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6788__A1 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout53_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5460__A1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _0454_ _0373_ _0460_ _0456_ _0465_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__4015__A2 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__I _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__I1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _0949_ _2631_ _2733_ _1646_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6960__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3958_ as2650.r0\[1\] _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6677_ _1498_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3889_ _3421_ _3423_ _3424_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6712__A1 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5515__A2 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ _1669_ _1673_ _1440_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5559_ _3306_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _0052_ clknet_leaf_53_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3829__A2 _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6779__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7293__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4254__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6481__C _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3677__I _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4006__A2 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7149__I _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5054__I1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6951__A1 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3765__A1 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5132__I _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4245__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ as2650.r0\[6\] as2650.r0\[5\] as2650.r0\[4\] as2650.r0\[3\] _1101_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5993__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4861_ _3173_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6600_ as2650.stack\[7\]\[10\] _2592_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3812_ _3326_ _3345_ _3347_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4792_ as2650.pc\[7\] _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6942__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3743_ _3152_ _3150_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6531_ _0471_ _2509_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3674_ as2650.ins_reg\[4\] _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6462_ _1128_ _1138_ _2472_ _2473_ _1504_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5413_ _1475_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6393_ _2303_ _2300_ _2376_ _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4181__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5344_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _0961_ _1369_ _1372_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7014_ _2983_ _2985_ _2987_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4226_ as2650.holding_reg\[5\] _0428_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4088_ _3410_ _0286_ _0292_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6630__B1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__I _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_37_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5984__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3995__A1 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5036__I1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5197__B1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3747__A1 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _3310_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__A1 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3960__I _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__S _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6492__B _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7100__C _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7189__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4966__I _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7101__A1 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__S _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4011_ _3539_ _3542_ _3544_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_77_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A3 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5415__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _0941_ as2650.pc\[1\] _0887_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3977__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7168__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5893_ _1765_ _1897_ _1904_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_90_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ _1013_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3729__A1 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4775_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5238__S _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6514_ _1537_ _2522_ _1633_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3726_ net10 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__A3 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _1004_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3657_ _3181_ _3192_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4154__A1 _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3588_ net53 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6376_ as2650.addr_buff\[0\] as2650.addr_buff\[1\] as2650.addr_buff\[2\] _2390_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5327_ _1403_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3780__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5258_ _0930_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4209_ _0287_ _3562_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5189_ _0676_ _0922_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4209__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5500__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7159__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6906__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5709__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6906__B2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__B _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4786__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5893__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6437__A3 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4448__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__B _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6373__A2 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _0667_ _0740_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4491_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6230_ _2129_ _2247_ _2127_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5884__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6161_ _1798_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7086__B1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5112_ as2650.stack\[4\]\[5\] _1230_ _1261_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6092_ _2111_ as2650.stack\[5\]\[4\] as2650.stack\[4\]\[4\] _2112_ _2113_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7204__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7354__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6994_ _2963_ _2969_ _2971_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6061__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5945_ _1968_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5876_ _1502_ _1317_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _3178_ _0850_ _0813_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5572__B1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _0939_ _0933_ _0940_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ _3149_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4689_ _0853_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6428_ _3237_ _3240_ _2439_ _3350_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _2372_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__A3 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4850__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4602__A2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4366__A1 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4118__A1 _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__C _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5405__I _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6815__B1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7377__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6291__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ _3487_ _3524_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5730_ _1760_ _1584_ _1763_ _1738_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _0874_ _1702_ _1703_ _3265_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7400_ _0223_ clknet_leaf_36_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4612_ _0707_ _0796_ _0797_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5592_ _0924_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7331_ _0154_ clknet_leaf_26_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ _0689_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7262_ _0085_ clknet_leaf_51_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4474_ _0625_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _2230_ _0473_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7193_ _0016_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _2110_ _2161_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6075_ _1125_ _1812_ _1007_ _1542_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5026_ _1160_ _0589_ _1194_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_113_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__B2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _0993_ _2636_ _2955_ _1939_ _2606_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_80_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__I _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5928_ _1662_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _1876_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4899__A2 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5934__B _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6749__C _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6273__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__B2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3626__A3 as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6025__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6576__A2 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__A1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__A1 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4354__A4 _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6659__C _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ _3400_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6264__A1 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6900_ _2206_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A1 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6831_ _2133_ _2766_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6567__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4578__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6762_ _2712_ _0312_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3974_ _3508_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ _1746_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6693_ _3267_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4214__I _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ _1683_ _1594_ _1684_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5575_ _1586_ _1617_ _1619_ _1621_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_89_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__C _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7314_ _0137_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4526_ _3362_ _0691_ _0716_ _0635_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _0068_ clknet_leaf_57_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4457_ _3159_ _0647_ _3229_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_132_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7176_ _1794_ _3124_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A4 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4388_ _0484_ _0487_ _0503_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3856__A3 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _0872_ _1740_ _2006_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6255__A1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _2040_ _2050_ _2079_ _2037_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _1161_ _1134_ _0540_ _0997_ _0490_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6007__A1 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4281__A3 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__C _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5230__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4124__I _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6730__A2 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6494__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6246__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7415__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__B _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3783__A2 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ as2650.cycle\[2\] _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6182__B1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _1428_ _0814_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _0429_ _0442_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ _0995_ _1376_ _1381_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7030_ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4242_ _0412_ _0436_ _0444_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6788__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _0489_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5212__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6745_ _1222_ _1634_ _2727_ _2732_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ _3490_ _3491_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6960__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4971__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _1300_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3888_ _3412_ _3253_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5627_ net25 _0911_ _1670_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6712__A2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4723__A1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _1515_ _1488_ _1489_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _0689_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5489_ _1542_ _1530_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6476__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _0051_ clknet_leaf_40_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7159_ _1720_ _3110_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6228__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__A3 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6400__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3765__A2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4962__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4789__I _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__C _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5413__I _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__I _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5569__B _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _3318_ _1030_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3811_ as2650.psl\[3\] _3346_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_127_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4791_ _0967_ _0956_ _0968_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ _1150_ _2526_ _2537_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3742_ _3277_ _3226_ _3153_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4953__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4699__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6155__B1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _1096_ _3362_ _1158_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3673_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5412_ _1475_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6392_ _1246_ _0539_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5343_ _0675_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__A1 as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5274_ as2650.stack\[0\]\[5\] _1370_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ net45 _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4225_ as2650.holding_reg\[5\] _0428_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_101_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5681__A2 _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4156_ _3543_ _0328_ _0358_ _3300_ _3298_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__6863__B _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4087_ _3430_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6630__A1 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5433__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6630__B2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4492__I0 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3995__A2 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5197__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5197__B2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _2712_ _0313_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__3747__A2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4944__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__B1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6659_ _2641_ _2644_ _2645_ _2648_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__B _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6697__A1 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6449__A1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5661__C _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6492__C _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3688__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__B _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5360__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7101__A2 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__I _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6860__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4010_ _3543_ _3503_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5415__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6612__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _1885_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3598__I _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4912_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__A2 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5892_ _1912_ _1916_ _1419_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7168__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4843_ _3259_ _3364_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4931__B _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6915__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3729__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6513_ _1123_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3725_ as2650.halted _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6679__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6444_ _3317_ _2455_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3656_ _3182_ _3185_ _3187_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__7283__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5762__B _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ as2650.addr_buff\[3\] _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5326_ as2650.r123\[3\]\[0\] _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5257_ _0895_ _1253_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6851__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4457__A3 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4208_ _0403_ _0408_ _0411_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5188_ _1315_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4892__I _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4139_ as2650.r0\[3\] _0314_ _0320_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6603__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4090__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5590__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4132__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4145__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__I _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7095__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6842__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5581__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _0673_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4136__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5074__S _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _1989_ _2171_ _2178_ _1994_ _2048_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3895__A1 _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7086__A1 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5111_ _1262_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _1211_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5042_ _0927_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ net41 _2970_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6061__A2 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _1464_ _1466_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5757__B _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4826_ as2650.psl\[6\] _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5021__B1 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ as2650.stack\[6\]\[1\] _0934_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5572__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__B2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5048__I _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ _3171_ _3243_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _3206_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3639_ _3174_ _3150_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6358_ _1246_ _2371_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5309_ _0961_ _1390_ _1393_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _2302_ _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A2 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7179__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4063__A1 _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6770__C _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4366__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5866__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__A1 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7068__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3629__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__B _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6291__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6043__A2 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _3487_ _3524_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5577__B _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _1675_ _1029_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ as2650.r123_2\[2\]\[7\] _0738_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5591_ net53 _1636_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7330_ _0153_ clknet_leaf_26_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _0725_ _0690_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7261_ _0084_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5306__A1 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _0663_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6212_ _1185_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5857__A2 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4500__I _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _0015_ clknet_leaf_66_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3868__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7059__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _1209_ as2650.stack\[3\]\[5\] as2650.stack\[2\]\[5\] _1920_ _2162_ _2163_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7321__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6806__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6074_ _1225_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__B _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5025_ _1169_ _1181_ _1193_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4832__A3 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _1249_ _2787_ _2954_ _1443_ _2410_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5793__A1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5927_ _1949_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4391__B _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _1833_ _1422_ _1596_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4809_ as2650.stack\[6\]\[9\] _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4348__A2 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _0447_ _1025_ _1026_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3859__A1 _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5241__I _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6025__A2 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3696__I _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4992__C1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7344__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5839__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__I _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _2806_ _2813_ _2814_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6761_ _1184_ _0361_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5775__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _3148_ _3365_ _3222_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6972__B1 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5712_ _3195_ _1488_ _3200_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6692_ _2641_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5527__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5643_ _3304_ _1416_ _1685_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5574_ _1620_ _1056_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7313_ _0136_ clknet_leaf_62_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4525_ _0365_ _0693_ _0714_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7244_ _0067_ clknet_leaf_51_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _3141_ _3170_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ as2650.psu\[0\] _3121_ _3123_ _3100_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ _2139_ _2144_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3856__A4 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _2049_ _2067_ _2077_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ as2650.psl\[5\] _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4018__A1 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5929__C _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7217__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6959_ _1247_ _2787_ _2938_ _2790_ _1887_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6620__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7367__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6191__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6776__B _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6494__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6246__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4257__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5057__I0 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5757__A1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6016__B _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4310_ _0433_ _0437_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ as2650.stack\[0\]\[12\] _1377_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4241_ _0271_ _0301_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__A2 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__S _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4172_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6788__A3 _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5996__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5996__B2 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6813_ _2693_ _2797_ _1847_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5748__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__B2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3956_ _3487_ _3489_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6744_ _1833_ _2047_ _2730_ _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _2628_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3887_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5626_ _1671_ _1442_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6173__A1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5557_ _1156_ _1601_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5056__I _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__B2 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ _3493_ _0690_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ as2650.addr_buff\[4\] _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6476__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4439_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7227_ _0050_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4487__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7158_ _3084_ _3105_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _1885_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4239__A1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7089_ _0418_ _0422_ _3041_ _3047_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6615__I _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6400__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4411__A1 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5675__B _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3974__I _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4962__A2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6164__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5911__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7130__B _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__I _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3810_ as2650.carry _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ as2650.stack\[6\]\[6\] _0957_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3741_ _3225_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6460_ _2465_ _3348_ _2468_ _2470_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6155__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3672_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6155__B2 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5411_ _1476_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6391_ _2332_ _2375_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5342_ _0928_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6458__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ _0954_ _1369_ _1371_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4469__A1 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7012_ _2968_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5130__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _0359_ _0328_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3692__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6863__C _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _0287_ _3273_ _3426_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6630__A2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__I1 as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5197__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _1041_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6727_ _2679_ _2713_ _2714_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3939_ _3463_ _3467_ _3436_ _3473_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4944__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _2647_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6146__B2 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6697__A2 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _1438_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _0961_ _2584_ _2587_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6449__A2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3969__I _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6385__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6137__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__A2 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3879__I _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__A2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _1889_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4623__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _1081_ _0868_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5891_ _1436_ _1914_ _1915_ _1517_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6376__A1 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _0812_ _0800_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5718__A4 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ as2650.pc\[4\] _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3724_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _1159_ _2520_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7428__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6679__A2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _3188_ _3190_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6443_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6374_ _2384_ _2387_ _1640_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4154__A3 _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5325_ _0994_ _1397_ _1402_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5256_ _0796_ _1351_ _1359_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ _0293_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6851__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4457__A4 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__S _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5187_ _0833_ _1304_ _1312_ _1130_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _3257_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3789__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6603__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4069_ _3399_ _3584_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4614__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6367__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5590__A2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5953__B _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7095__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4853__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3656__A2 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__A1 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5581__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6530__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ as2650.stack\[4\]\[4\] _1226_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _1251_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6694__B _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5090__S _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4844__A1 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _2968_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5943_ _1940_ _1964_ _1966_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6349__A1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5874_ _1108_ _1442_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7010__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7250__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4825_ _0995_ _0982_ _0996_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5021__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5021__B2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5572__A2 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3707_ _3217_ _3231_ _3242_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4687_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3638_ as2650.cycle\[1\] _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6426_ _0655_ _0637_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5324__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6357_ _0985_ _2330_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__A2 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ as2650.stack\[1\]\[5\] _1391_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _2303_ _2259_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6824__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _1349_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4835__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4063__A2 _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4143__I _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6760__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6512__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5946__S0 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3877__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__B1 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3629__A2 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__C _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7273__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5858__B _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4610_ _0577_ _0627_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5590_ _1566_ _0907_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5554__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ _0726_ _0727_ _0730_ _0698_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4988__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7260_ _0083_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4472_ _3303_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6503__A1 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6211_ _2220_ _2222_ _2228_ _1707_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7191_ _0014_ clknet_leaf_66_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3868__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _1467_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A2 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _0948_ _2051_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _3134_ _0801_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4293__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ _2420_ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5093__I1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6443__I _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ as2650.pc\[1\] net6 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5793__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6990__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5857_ _1619_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _0931_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5545__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6742__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5788_ _1795_ _0904_ _1796_ _1819_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4739_ _0640_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _2420_ _2421_ _1639_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7389_ _0212_ clknet_leaf_44_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6618__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5522__I _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7296__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A2 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4992__B1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4992__C2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4802__S _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6760_ _1540_ _2684_ _0318_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6972__A1 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3972_ _3506_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5775__A2 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6972__B2 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5711_ _1738_ _3201_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6691_ _3570_ _3545_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5642_ _1014_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5573_ _1502_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5607__I _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4511__I _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7312_ _0135_ clknet_leaf_61_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4524_ _0656_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7243_ _0066_ clknet_leaf_51_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4455_ _3128_ _3132_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6866__C _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7174_ _1698_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4386_ net3 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6125_ _2141_ _2143_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5342__I _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6056_ _2033_ _2040_ _2034_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ _1170_ _3569_ _0376_ _3335_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A2 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _2382_ _2937_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _1208_ _1010_ _1926_ _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6889_ _2869_ _2871_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6715__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6715__B2 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6479__B1 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7140__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5454__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5057__I1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7311__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5509__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6182__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4193__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ _3410_ _0439_ _0443_ _0293_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5693__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6258__I _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4171_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4248__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5445__A1 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6812_ net34 _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4506__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5748__A2 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _1414_ _2402_ _0839_ _1222_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3955_ _3487_ _3489_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _2638_ _2660_ _2662_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3886_ _3368_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4971__A3 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _1000_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5556_ _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5781__B _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4507_ _3438_ _0691_ _0697_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7122__A1 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5487_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7226_ _0049_ clknet_leaf_40_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4438_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5684__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7157_ _3084_ _3085_ _3102_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4369_ _0403_ _0566_ _0570_ _0293_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6108_ _0955_ _1983_ _2128_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6228__A3 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7088_ _0299_ _0306_ _3042_ _3045_ _3046_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4239__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _3140_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3998__A1 _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7334__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6936__A1 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4962__A3 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6164__A2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4151__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4175__B2 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5911__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7113__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3989__A1 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6027__B _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4326__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3740_ _3266_ _3267_ _3273_ _3275_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6155__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3671_ as2650.ins_reg\[3\] _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5410_ _0669_ as2650.r123_2\[0\]\[0\] _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6390_ _1562_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _1410_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7104__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__S _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ as2650.stack\[0\]\[4\] _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7207__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4469__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7011_ _0363_ _2976_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ _0367_ _0370_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4154_ _3295_ _3359_ _3501_ _0282_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3692__A3 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7357__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4085_ _3272_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4236__I as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__A1 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6451__I _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _1533_ _3539_ _3542_ _3544_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3938_ _3409_ _3470_ _3472_ _3429_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6657_ _1746_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6146__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3869_ _3332_ _3131_ _3289_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5608_ _1653_ _1555_ _1595_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6588_ as2650.stack\[7\]\[5\] _2585_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3904__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5539_ _1034_ _1013_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7209_ _0032_ clknet_leaf_47_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6626__I _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5530__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A1 _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4148__A1 _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5705__I _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5648__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__A3 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__A2 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5890_ _1907_ _1908_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ _3178_ _0642_ _0807_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6376__A2 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__I _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ _0951_ _0933_ _0952_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _2516_ _0482_ _2519_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3723_ _3252_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6128__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4139__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6442_ _2437_ _2442_ _2453_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3654_ _3189_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6373_ _1767_ _2372_ _2386_ _2009_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4154__A4 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5324_ as2650.stack\[1\]\[12\] _1398_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5639__A1 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ as2650.r123_2\[1\]\[7\] _1354_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4206_ _0409_ _0330_ _0410_ _0403_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _0826_ _1304_ _1312_ _1314_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A2 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6446__I _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _3517_ _0321_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6064__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4068_ _0270_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4378__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _2631_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5953__C _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4302__A1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4853__A2 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5260__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4161__S0 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5581__A3 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__C _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4541__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6294__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _0893_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4844__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5170__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6046__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6046__B2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6991_ _2968_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _1318_ _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5873_ _0888_ _3373_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5006__C1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ as2650.stack\[6\]\[12\] _0983_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5021__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3706_ _3147_ _3238_ _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4686_ _0490_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6425_ _2436_ _1593_ _1602_ _1606_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3637_ _3155_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5345__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6356_ _2366_ _2369_ _0867_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _0954_ _1390_ _1392_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6287_ as2650.pc\[8\] _2230_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5238_ _0669_ as2650.r123_2\[1\]\[0\] _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5627__A4 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6176__I _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4063__A3 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6760__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_30_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__S1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__A1 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7418__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5858__C _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5787__B1 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6200__A1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6751__A2 _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4540_ _0482_ _0644_ _0729_ _0657_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4471_ _3206_ _0649_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5165__I _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6503__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ _2225_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4514__A1 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7190_ _0013_ clknet_leaf_66_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _2111_ as2650.stack\[1\]\[5\] as2650.stack\[0\]\[5\] _0929_ _2161_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5314__I0 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _1988_ _2092_ _1996_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5023_ _0315_ _0261_ _1002_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6019__A1 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6724__I _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6974_ _1740_ _2944_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5242__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ as2650.pc\[0\] net5 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6990__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4244__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _3246_ _1024_ _1037_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _0932_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5787_ _1800_ _1815_ _1817_ _1818_ _1571_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4738_ _3207_ _0918_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _0378_ _1424_ _1671_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7388_ _0211_ clknet_leaf_44_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _2239_ _2352_ _2353_ _2162_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4419__I _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6430__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5784__A3 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A1 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4992__B2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6497__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6972__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7390__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6421__A1 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6421__B2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3971_ _3505_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6972__A2 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4064__I _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ _0874_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4983__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6690_ _1172_ _3525_ _3526_ _2642_ _2643_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _3260_ _1516_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6185__B1 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4735__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _0806_ _0852_ _1500_ _1618_ as2650.halted _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_117_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7311_ _0134_ clknet_leaf_64_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4523_ _3567_ _0694_ _0644_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4013__B _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7242_ _0065_ clknet_leaf_53_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4454_ _3250_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__A1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6719__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _1305_ _3104_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ _3325_ _3423_ _3347_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_98_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6124_ _2141_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _0866_ _2071_ _2076_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6660__A1 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ as2650.psl\[1\] _1173_ _1174_ _3325_ _3432_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__5779__B _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A3 _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _1740_ _2926_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6963__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4974__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5908_ _1927_ _1932_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6888_ _2275_ _2870_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5839_ _0826_ _1157_ _1708_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4726__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__B1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6479__A1 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6479__B2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7263__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7140__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3701__A2 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5454__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6403__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5206__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3937__B _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__B1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4717__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4193__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__A2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7144__B _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6890__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__B2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ net9 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6642__A1 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5445__A2 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6811_ net51 _2739_ _2740_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4956__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _1040_ _2402_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3954_ _3416_ _3386_ _3488_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_108_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6673_ _2661_ _1950_ _1788_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3885_ _3255_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5618__I _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ _0910_ _0925_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7286__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5555_ _1080_ _1578_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4506_ _0633_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3931__A2 _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5486_ _1184_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7122__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _0048_ clknet_leaf_40_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4437_ _3237_ _3240_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4487__A3 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7156_ _3083_ _3108_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4368_ _3410_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _1984_ _2126_ _2127_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7087_ _0277_ _3044_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _0501_ _0481_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6633__A1 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6038_ _2005_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3601__I _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6117__C _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4962__A4 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3922__A2 _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7113__A2 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6359__I _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5675__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3686__A1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6624__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6094__I _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3989__A2 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6027__C _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7139__B _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ _3194_ _3202_ _3205_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_118_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6978__B _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ as2650.r123\[3\]\[7\] _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7104__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ _1361_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ _2972_ _0472_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6863__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4222_ _0356_ _0424_ _0426_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4153_ _0357_ _0327_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6218__B _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__A1 _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4986_ _0589_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6725_ _3539_ _3542_ _3544_ _1533_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3937_ _3255_ _3361_ _3409_ _3471_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4252__I _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6656_ _0317_ _1605_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3868_ _3316_ _3145_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_137_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__B _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5607_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _0954_ _2584_ _2586_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3799_ _3329_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _0850_ _1553_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_121_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _1525_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7208_ _0031_ clknet_leaf_45_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _3091_ _3093_ _1794_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7301__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4148__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6089__I _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5721__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4337__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__A2 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5820__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4840_ _3194_ _3158_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6376__A3 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ as2650.stack\[6\]\[3\] _0934_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5584__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6510_ _1098_ _0726_ _2517_ _2518_ _1121_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3722_ _3141_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6441_ _2444_ _2448_ _2451_ _2452_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_88_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3653_ as2650.ins_reg\[7\] _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4800__I _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6372_ _0989_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3898__A1 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7089__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5323_ _0990_ _1397_ _1401_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7324__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6836__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5639__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5254_ _1358_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4205_ _0396_ _3421_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4311__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ _1313_ _1307_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4136_ _3376_ _0330_ _0341_ _3168_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6064__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ _0271_ _0272_ _0273_ _3480_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _1124_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6708_ _2498_ _1579_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _2610_ _2621_ _2629_ _1204_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4550__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6827__A1 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4302__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4157__I _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5697__B _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4161__S1 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3813__A1 _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6366__I0 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7347__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__A3 _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A2 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__A1 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6990_ _1561_ _2437_ _2966_ _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_93_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _1609_ _1951_ _1943_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3804__A1 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5872_ _1640_ _1891_ _1894_ _1896_ _0890_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__5006__B1 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4823_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5557__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4754_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3705_ _3240_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5309__A1 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4685_ as2650.r0\[5\] _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _1081_ _0838_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3636_ _3147_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6355_ _1458_ _2367_ _2368_ _1469_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6809__A1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ as2650.stack\[1\]\[4\] _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6286_ _2300_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5237_ _1347_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6457__I _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4296__A1 as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5168_ _0640_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4119_ as2650.r123\[0\]\[4\] as2650.r123\[2\]\[4\] as2650.r123_2\[0\]\[4\] as2650.r123_2\[2\]\[4\]
+ _3143_ _3137_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _1253_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5548__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5536__I _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5980__B _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5271__I _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4287__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5787__B2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4615__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5539__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4211__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__B net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _3391_ _0632_ _0661_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6986__B _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5711__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ as2650.stack\[7\]\[5\] as2650.stack\[4\]\[5\] as2650.stack\[5\]\[5\] as2650.stack\[6\]\[5\]
+ _1972_ _2111_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6267__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6071_ _1902_ _2084_ _2091_ _1994_ _1753_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5022_ as2650.psu\[0\] _1175_ _0760_ as2650.psu\[5\] _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4953__C _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _1600_ _2948_ _2951_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _0810_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__A1 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5855_ _1878_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5786_ _1603_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _3281_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5356__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4668_ _0821_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3619_ _3153_ _3154_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ as2650.addr_buff\[4\] _1945_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5702__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7387_ _0210_ clknet_leaf_43_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4599_ _0530_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3805__S _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ as2650.stack\[7\]\[10\] _2115_ _1920_ as2650.stack\[6\]\[10\] _2353_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6269_ _1457_ _2285_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3604__I _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5959__C _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7192__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A2 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6650__I _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4170__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ net6 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4432__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4983__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6185__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _0913_ _0908_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6185__B2 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _1032_ _1045_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4735__A2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7310_ _0133_ clknet_leaf_61_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4522_ _0711_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4453_ _3182_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7241_ _0064_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ _1305_ _1643_ _3102_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4384_ _0481_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6123_ _0759_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _1210_ as2650.stack\[3\]\[3\] as2650.stack\[2\]\[3\] _1930_ _2075_ _2076_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_100_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _3372_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6660__A2 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6412__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6956_ _2211_ _2378_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5907_ _1921_ _1928_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4974__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6887_ _2866_ _2868_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ as2650.psu\[7\] _1157_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5923__A1 _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__B2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _1551_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6479__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6100__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6645__I _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4593__C _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6167__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6167__B2 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4717__A2 _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7131__A3 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5142__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A3 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4653__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4075__I _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6810_ _2635_ _2793_ _2795_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6741_ _1174_ _1801_ _2728_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3953_ _3385_ _3234_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4956__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6672_ _2661_ _1950_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3884_ _3347_ _3419_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5623_ _1156_ _1318_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5554_ _1515_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _0321_ _0693_ _0696_ _0657_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5485_ _1537_ _1524_ _1539_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7122__A3 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4436_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7224_ _0047_ clknet_leaf_43_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7155_ as2650.psu\[4\] _3103_ _3107_ _3096_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ as2650.holding_reg\[7\] _3273_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3695__A2 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _0883_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ _3455_ _1086_ _0277_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ as2650.holding_reg\[6\] _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__B _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6633__A2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _1908_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6397__A1 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _1244_ _2665_ _2919_ _2623_ _1582_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7230__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5972__C _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7380__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4883__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3686__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3999__I _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4635__A1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5719__I _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6560__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _1362_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6312__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6312__B2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4221_ as2650.r123\[2\]\[4\] _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6863__A2 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ _3368_ _3458_ _3532_ _3560_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_110_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3702__I _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4626__A1 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6218__C _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7253__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4929__A2 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _0773_ _1144_ _1153_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6724_ _0336_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3936_ _3460_ _3255_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6655_ _3507_ _2640_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3867_ _3402_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5606_ _1097_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6551__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ as2650.stack\[7\]\[4\] _2585_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3798_ _3329_ as2650.r123_2\[0\]\[7\] _3330_ _3333_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7065__B _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5537_ _3365_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5364__I _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5468_ _1522_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6303__B2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7207_ _0030_ clknet_leaf_47_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6854__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4419_ _0609_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5399_ _0896_ _0927_ as2650.stack_ptr\[2\] _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7138_ _1710_ _3077_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__B _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4708__I _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7069_ _0870_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5032__C _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A2 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7031__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4443__I _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4856__A1 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4608__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7276__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5820__A3 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5033__B2 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5584__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _3245_ _3247_ _3251_ _3256_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6440_ _1034_ _1021_ _1038_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3652_ as2650.ins_reg\[6\] _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6533__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _1243_ _2344_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5184__I _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3898__A2 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7089__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ as2650.stack\[1\]\[11\] _1398_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6836__A2 _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5639__A3 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5253_ _0783_ as2650.r123_2\[1\]\[6\] _1348_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__A1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ _3421_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5184_ _1129_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _3352_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4066_ _3582_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5787__C _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5024__A1 _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6772__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4968_ _1127_ _1133_ _1137_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6707_ _1600_ _2690_ _2692_ _2693_ _2695_ _1847_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_71_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3919_ as2650.holding_reg\[1\] _3269_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4899_ _0560_ _3345_ _0569_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _2623_ _2627_ _2628_ _0890_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6524__A1 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3607__I _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _1141_ _2463_ _1665_ _0591_ _2573_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__3889__A2 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__A2 _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5822__I _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7299__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5263__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3813__A2 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__A2 _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4173__I _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5318__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__I1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6515__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6049__B _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5940_ _1639_ _1944_ _1954_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_94_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5179__I _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4083__I _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__B2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4822_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4753_ as2650.pc\[1\] _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4811__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ as2650.addr_buff\[7\] _3239_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6506__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4684_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _0994_ _1886_ _2435_ _1695_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3635_ _3170_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6354_ as2650.stack\[7\]\[11\] _2115_ _2195_ as2650.stack\[6\]\[11\] _2368_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3740__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _1382_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6285_ _0979_ _1186_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5236_ _0672_ _0682_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5493__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _3180_ _0917_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ _3127_ _0322_ _0323_ _3131_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5098_ _1210_ _0930_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5245__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4049_ _3581_ _3582_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6406__C _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__A1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5548__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7170__A1 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7170__B2 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5720__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6648__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5484__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4168__I _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5236__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4039__A2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3800__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5787__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5539__A2 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5727__I _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4631__I _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7161__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5663__S _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A2 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6070_ _2086_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5021_ _1182_ _1134_ _3569_ _1183_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5078__I1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__I _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _2814_ _2944_ _2950_ _1821_ _2479_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3710__I _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6975__A1 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5923_ _3507_ _1945_ _1946_ _1528_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5854_ _1042_ _1033_ _1019_ _1797_ _1306_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4805_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5637__I _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5785_ _1029_ _1816_ _1805_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4736_ _0912_ _0915_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_119_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4667_ _0850_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6406_ _2053_ _2409_ _2418_ _1052_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3618_ as2650.cycle\[3\] as2650.cycle\[2\] _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7386_ _0209_ clknet_leaf_47_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4598_ _0784_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7073__B _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6337_ _2199_ as2650.stack\[5\]\[10\] as2650.stack\[4\]\[10\] _1252_ _2352_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__I _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6268_ _1972_ as2650.stack\[5\]\[8\] as2650.stack\[4\]\[8\] _0897_ _2285_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _0962_ _1334_ _1337_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ _2211_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4716__I _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6718__B2 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__I _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5941__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3704__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5282__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5209__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4680__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4432__A2 _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__A3 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6185__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ _1445_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ _0650_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7134__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7240_ _0063_ clknet_leaf_42_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4452_ _3183_ _3186_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _1794_ _3120_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3705__I _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4383_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5192__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _3140_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A1 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _2023_ _2073_ _2074_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5999__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _0336_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4120__A1 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4671__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4536__I _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _1414_ _1296_ _2609_ _2934_ _1755_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5620__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _0894_ as2650.stack\[3\]\[0\] as2650.stack\[2\]\[0\] _1930_ _1469_ _1931_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6886_ _2274_ _2866_ _2868_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7068__B _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5837_ _1861_ _1862_ net4 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5367__I _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5923__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3934__A1 _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4719_ _3198_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7125__A1 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5699_ _1712_ _1733_ _1734_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7369_ _0192_ clknet_leaf_39_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3615__I _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5439__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5830__I _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6939__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6939__B2 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__B _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4414__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4178__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7116__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4102__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A4 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5602__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__A2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _1739_ _2711_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3952_ _3486_ _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4956__A3 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6671_ as2650.pc\[0\] net5 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6158__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3883_ _3414_ _3418_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5622_ _1651_ _1667_ net25 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5553_ _1490_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7107__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__I _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4504_ _3514_ _0694_ _0692_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5484_ _1538_ _1530_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7223_ _0046_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4435_ _3335_ _3263_ _3146_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_104_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7182__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4341__A1 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7154_ _1723_ _3106_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4366_ _3272_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4975__B _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3695__A3 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6105_ _2084_ _2093_ _2125_ _2037_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _1022_ _3504_ _3043_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4297_ _0356_ _0499_ _0500_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7070__C _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6036_ _1894_ _2052_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5841__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4266__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6397__A2 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _2666_ _2337_ _2918_ _2626_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _2705_ _2852_ _2826_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5097__I _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3907__A1 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6430__B _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4580__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4885__B _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5832__A1 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4635__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4399__A1 _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5899__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5899__B2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7104__A4 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4323__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4220_ _3450_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4874__A2 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4151_ _3286_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6076__A1 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _0282_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4626__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6379__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4929__A3 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4984_ _1004_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6723_ _2707_ _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3935_ _3464_ _3469_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ _2642_ _2643_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3866_ _3401_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _1445_ _1630_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6250__B _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6585_ _2576_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5645__I _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3797_ _3332_ _3132_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6551__A2 _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5536_ _1552_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7065__C _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5467_ as2650.addr_buff\[0\] _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4314__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7206_ _0029_ clknet_leaf_46_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4418_ _0607_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _1464_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3912__I1 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7137_ _0798_ _0878_ _1709_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _3315_ _0535_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6067__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7068_ _0873_ _3014_ _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _3247_ _1299_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6790__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_64_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4553__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4305__A1 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__A2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5105__I0 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5805__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4608__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4634__I _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3720_ _3252_ _3255_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5893__C _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3651_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5465__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _1810_ _2380_ _2383_ _0822_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5321_ _0986_ _1397_ _1400_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _0770_ _1351_ _1357_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5639__A4 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4847__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ _0401_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5183_ _1165_ _1304_ _1308_ _1312_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _3366_ _0334_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4065_ _3580_ _3535_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5009__C1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4967_ _1041_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6772__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6706_ _1990_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3918_ _3283_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4898_ _1066_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6637_ _2266_ _1427_ _2622_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3849_ as2650.addr_buff\[5\] _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6524__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _1157_ _1138_ _1202_ _2572_ _1504_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_118_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ _1567_ _1568_ _1518_ _1565_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6499_ _0725_ _2455_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__A2 _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3623__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3821__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4526__A1 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A1 _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__B2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7243__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4629__I _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6844__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7393__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _1441_ _0925_ _1767_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4821_ as2650.pc\[12\] _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6754__A2 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4752_ _0892_ _0933_ _0935_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4765__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3703_ as2650.cycle\[7\] _3196_ _3200_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5195__I _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4683_ _0636_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6506__A2 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6422_ _1888_ _2401_ _2434_ _1981_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3634_ _3135_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6353_ _0929_ as2650.stack\[5\]\[11\] as2650.stack\[4\]\[11\] _0898_ _2367_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5304_ _1383_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3740__A2 _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ _1240_ _2230_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5235_ _0995_ _1341_ _1346_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5166_ _1032_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4117_ as2650.r0\[4\] _3332_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5097_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6442__A1 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ as2650.holding_reg\[2\] _3533_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ as2650.stack\[7\]\[2\] _1465_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5548__A3 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6422__C _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4508__A1 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7266__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5181__A1 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__A1 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__B2 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4119__S0 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5236__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6984__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6736__A2 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4380__C1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _1188_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6574__I _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6971_ _2408_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4308__B _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5922_ _1498_ _1051_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5853_ _3214_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ as2650.pc\[9\] _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4738__A1 _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4822__I _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5784_ _1022_ _3318_ _1144_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7289__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _3181_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_120_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _0621_ _0837_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _2264_ _2400_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3617_ as2650.cycle\[7\] as2650.cycle\[6\] as2650.cycle\[5\] as2650.cycle\[4\] _3153_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_128_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7385_ _0208_ clknet_leaf_58_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5653__I _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4597_ _0783_ as2650.r123_2\[2\]\[6\] _0684_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6336_ _1782_ _2346_ _2350_ _1779_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ as2650.stack\[7\]\[8\] _1465_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5218_ as2650.stack\[2\]\[5\] _1335_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6198_ _2212_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6484__I _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ as2650.stack\[3\]\[6\] _1283_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3901__I _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5218__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6415__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__A1 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6718__A2 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5828__I _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7143__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6406__A1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5209__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6957__A2 _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7431__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3640__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _3570_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5473__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6893__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7170_ as2650.psu\[1\] _3117_ _3119_ _3100_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4382_ as2650.r0\[7\] _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6121_ _2103_ _2105_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _1968_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__I _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4120__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6948__A2 _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6954_ _2375_ _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4980__C _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5620__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5905_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6253__B _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6885_ _2652_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4552__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5836_ _1719_ _1003_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4187__A2 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4718_ _3151_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5698_ _0560_ _1712_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7125__A2 _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6700__C _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7437_ _0260_ clknet_leaf_22_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4649_ _3187_ _0812_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6884__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7368_ _0191_ clknet_leaf_38_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6319_ _2303_ _2300_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7299_ _0122_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7304__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6636__B2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6939__A2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3870__A1 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7061__A1 _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4462__I _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7116__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5507__B _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__D _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6627__A1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4637__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4102__A2 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5850__A2 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5669__S _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A1 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ _3295_ _3359_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5468__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6670_ _2612_ _2639_ _2657_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ _3415_ _3416_ _3417_ _3413_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1654_ _1625_ _1661_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5366__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3916__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5552_ _0315_ _0817_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4503_ _3506_ _0651_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ as2650.addr_buff\[3\] _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7327__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6866__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4434_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7222_ _0045_ clknet_leaf_43_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7153_ _3072_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4365_ _0556_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _2092_ _2109_ _2124_ _1850_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ _3580_ _1022_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ as2650.r123\[2\]\[5\] _0425_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _2055_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5841__A2 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _1535_ _2139_ _2917_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _1646_ _2848_ _2850_ _2250_ _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4215__C _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ _1601_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6711__B _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _2769_ _2781_ _2784_ _2638_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3907__A2 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6306__B1 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6857__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6609__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4096__B2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__A1 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4399__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4141__B _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _3287_ _0354_ _0355_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6076__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4081_ as2650.holding_reg\[3\] _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5123__I1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3834__A1 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__I _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _0584_ _1093_ _1027_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ net30 net52 net28 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3934_ _3347_ _3468_ _3414_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6653_ _1171_ _3486_ _3524_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_3865_ _3220_ _3191_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5604_ _1149_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4011__A1 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _3331_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6584_ _2577_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6250__C _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _1582_ _1035_ _0852_ _1556_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5466_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4417_ _0354_ _0608_ _0614_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7205_ _0028_ clknet_leaf_57_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5511__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _1272_ _1454_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7136_ _1064_ _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4348_ _3313_ _0546_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6067__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4277__I _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7067_ _1012_ _3020_ _3021_ _3026_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5114__I1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4279_ _0332_ _3561_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _0947_ _1985_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7016__A1 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5610__B _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5578__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4740__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__A1 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6160__C _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4553__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__A1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5750__B2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4305__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5502__A1 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4388__S _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__A3 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__I1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4069__A1 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A2 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7007__A1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5018__B1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5569__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4241__A1 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5746__I _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__I _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3650_ as2650.ins_reg\[5\] _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5741__A1 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5741__B2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5682__S _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5320_ as2650.stack\[1\]\[10\] _1398_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6297__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ as2650.r123_2\[1\]\[5\] _1354_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4202_ _0263_ _0404_ _0405_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_87_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6049__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4133_ _0338_ _3366_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ _3478_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4480__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__B1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__I0 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6705_ _1991_ _2662_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3917_ _3287_ _3448_ _3452_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6261__B _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _0404_ _1067_ _0405_ _0406_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_71_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _2402_ _1898_ _2624_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3848_ _3317_ _3322_ _3381_ _3383_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5732__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3779_ _3312_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6567_ _1182_ _0848_ _2571_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ _1052_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6498_ _1650_ _2492_ _2507_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5449_ _3264_ _1502_ _1503_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__4299__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _1642_ _0829_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5799__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7195__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__A2 _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4820_ _0991_ _0982_ _0992_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ as2650.stack\[6\]\[0\] _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5962__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__I _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3702_ _3237_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4682_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ _3168_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6421_ _2411_ _2425_ _2433_ _1453_ _1939_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5714__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6352_ _1458_ _2364_ _2365_ _2159_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5303_ _0950_ _1384_ _1389_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6283_ _1240_ _2298_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3740__A3 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3724__I _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ as2650.stack\[2\]\[12\] _1342_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _3151_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ as2650.r123\[1\]\[4\] as2650.r123_2\[1\]\[4\] _3137_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4047_ _3580_ _3533_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5253__I0 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5998_ _1998_ _2007_ _2008_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5548__A4 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5953__A1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _0462_ _0785_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6619_ _2609_ _1898_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3634__I _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__I _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6130__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__A2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4119__S1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6613__C _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3809__I _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7210__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4380__C2 _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6970_ _2404_ _2913_ _2406_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__A1 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5921_ _1558_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ _1165_ _0845_ _0828_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6188__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6188__B2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _0978_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4738__A2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3719__I _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _1573_ _1808_ _1809_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4734_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _3181_ _3211_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6404_ as2650.addr_buff\[4\] _2416_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3616_ as2650.cycle\[1\] _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7384_ _0207_ clknet_leaf_56_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6360__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _0781_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6335_ _2006_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _1655_ _2273_ _2282_ _1940_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5217_ _0955_ _1334_ _1336_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6197_ _2213_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _0962_ _1282_ _1285_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4285__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ _1239_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6179__B2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__S _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7233__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7383__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A3 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6351__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__B2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6103__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6675__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4665__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6406__A2 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4417__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4923__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4432__A4 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5754__I _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4450_ _3158_ _0642_ _0628_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6342__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6893__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4381_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6120_ _0375_ _2104_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6585__I _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2072_ as2650.stack\[1\]\[3\] as2650.stack\[0\]\[3\] _1212_ _2073_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4656__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__A1 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__CLK clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _2333_ _2914_ _2376_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ _1919_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5620__A3 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6884_ _1135_ _0600_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3631__A2 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5908__A1 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5835_ _0853_ _0831_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6581__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4717_ _3174_ _3278_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5697_ _1324_ _1714_ _1199_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _0259_ clknet_leaf_20_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5136__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6884__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ _0190_ clknet_leaf_38_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4579_ _0719_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4895__A1 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7298_ _0121_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6636__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6249_ _0817_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5105__S _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__I0 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6428__C _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3870__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_58_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7061__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4743__I as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__B _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6324__A1 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5686__I0 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7279__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4139__B _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A3 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ _3283_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3881_ _3407_ _3269_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5620_ _1663_ _0819_ _1664_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_108_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5551_ _1301_ _1500_ _1518_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _0652_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5482_ _1174_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7221_ _0044_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6866__A2 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4433_ _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7152_ _3104_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4364_ _0557_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6103_ _2033_ _2084_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _3455_ _3483_ _3439_ _3445_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4295_ _3453_ _0453_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6034_ _1132_ _1499_ _1946_ _1538_ _1620_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3852__A2 _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6936_ _2667_ _2903_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6867_ _1235_ _2636_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6003__B1 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5818_ _1842_ _1844_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6798_ _2611_ _2783_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7095__B _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__B _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5394__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5749_ _1438_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7419_ _0242_ clknet_leaf_1_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4868__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7421__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3642__I _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__A2 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6793__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__A2 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3753__S _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__I _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4080_ _0284_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A3 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3834__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5479__I as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4383__I _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6784__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _1063_ _1085_ _1077_ _0854_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _2042_ _2708_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3933_ _3254_ _3368_ _3424_ _3408_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_3_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _3371_ _3302_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3864_ _3399_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6536__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _1632_ _1648_ _1649_ _1473_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6583_ _0950_ _2578_ _2583_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4011__A2 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3795_ _3125_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5534_ _1143_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7204_ _0027_ clknet_leaf_57_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4416_ as2650.r123\[1\]\[3\] _0610_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4314__A3 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5511__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ _1462_ _1458_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7135_ _1313_ _3085_ _3077_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4347_ _3393_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ _3022_ _3024_ _3025_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4278_ _0457_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5275__A1 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6017_ _0945_ _1983_ _2039_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6775__B2 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ net37 _2607_ _1151_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6527__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__D _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4002__A2 _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__A4 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4069__A2 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5520__C _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5018__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5018__B2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7317__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6766__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5569__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4241__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5741__A2 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5250_ _0754_ _1350_ _1356_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _0273_ _0266_ _0283_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_142_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5181_ _1303_ _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _3478_ _3479_ _3397_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6526__C _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5009__B2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4480__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__I _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6542__B _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6704_ _2611_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3916_ as2650.r123\[2\]\[0\] _3451_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4896_ _3418_ _3464_ _0262_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3847_ _3382_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1160_ _2469_ _0808_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3778_ _3313_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5732__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__I _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6497_ _2497_ _2499_ _2506_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5448_ _0315_ _0318_ _1299_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5496__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5379_ _1444_ _1445_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7118_ _1002_ _0831_ _1056_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5248__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7049_ _3171_ _1307_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5799__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6996__A1 _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7173__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4198__I _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__B _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4926__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6987__A1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__B1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6739__A1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _0931_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5962__A2 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3701_ _3232_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3973__A1 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7164__A1 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _3161_ _0811_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6420_ _0867_ _2401_ _2432_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3632_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5714__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _0894_ as2650.stack\[3\]\[11\] as2650.stack\[2\]\[11\] _2195_ _2365_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5302_ as2650.stack\[1\]\[3\] _1385_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6282_ _0974_ _2251_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3740__A4 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5233_ _0991_ _1341_ _1345_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4150__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _0995_ _1289_ _1294_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ _3535_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6978__A1 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5095_ _0896_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ as2650.holding_reg\[2\] _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6442__A3 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4453__A2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _1297_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4571__I _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4948_ _0773_ _1118_ _0321_ _3562_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__5953__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7155__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4879_ _1044_ _1046_ _1047_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7155__B2 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _1742_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6549_ _2510_ _2553_ _2554_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5469__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4141__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3650__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5641__A1 _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__A3 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6910__B _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3825__I _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4380__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4435__A2 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ _1892_ _1942_ _1943_ _1893_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _1688_ _1871_ _1872_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__5487__I _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ _0977_ as2650.stack\[6\]\[8\] _0932_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _1811_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3946__A1 _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4733_ _3133_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7137__A1 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _0843_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6403_ _2389_ _2279_ _2390_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3615_ _3150_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7383_ _0206_ clknet_leaf_56_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4595_ _0528_ _0667_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6360__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6334_ as2650.addr_buff\[2\] _2348_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4371__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _2280_ _2281_ _2060_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ as2650.stack\[2\]\[4\] _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6196_ _2173_ _2177_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4674__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5147_ as2650.stack\[3\]\[5\] _1283_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ as2650.stack\[5\]\[8\] _1237_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5623__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4029_ _3366_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5926__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__A1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6730__B _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7143__A4 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3645__I _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4362__A1 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4901__A3 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__I _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A2 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5614__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5100__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5917__A2 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3928__A1 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7119__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6590__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ _0556_ _0454_ _0579_ _0456_ _0581_ _3300_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_98_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4105__A1 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5153__I0 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6050_ _0896_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6087__B _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _3505_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4386__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5853__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4656__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6952_ _1605_ _2926_ _2931_ _2638_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5903_ _1253_ as2650.stack\[1\]\[0\] as2650.stack\[0\]\[0\] _1411_ _1928_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6883_ _2807_ _2810_ _2865_ _2841_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_81_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5620__A4 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3631__A3 _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5834_ _1795_ _3306_ _1796_ _1860_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5908__A2 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6030__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5765_ _3185_ _1577_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6550__B _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4592__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ _0678_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5696_ _1732_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7435_ _0258_ clknet_3_2_0_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _0677_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4344__A1 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _0189_ clknet_leaf_38_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4578_ _0471_ _0710_ _0632_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6317_ _0985_ _0538_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7297_ _0120_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6097__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6097__B2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6248_ _2264_ _2261_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5695__I1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _0894_ as2650.stack\[3\]\[6\] as2650.stack\[2\]\[6\] _2195_ _2197_ _2198_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7200__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5121__S _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7350__CLK clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6021__A1 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6572__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4583__A1 as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6088__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5686__I1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4934__I _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3880_ _3294_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A1 _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__A1 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _1593_ _1594_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _1534_ _1524_ _1536_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6315__A2 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _0043_ clknet_leaf_59_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4432_ _3141_ _3265_ _3276_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5714__B _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6596__I _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7151_ _0876_ _0877_ _1707_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4363_ _0505_ _0515_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6079__A1 _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _2114_ _2117_ _2121_ _2122_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6529__C _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7082_ _0299_ _0306_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _3314_ _0467_ _0497_ _3485_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7223__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5826__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _2053_ _2046_ _2054_ _1433_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5005__I _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7373__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6935_ _2904_ _2912_ _2915_ _1857_ _2457_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _1235_ _2787_ _2849_ _2790_ _2217_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_74_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6003__B2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5817_ _1842_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6797_ net51 _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6554__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ _1779_ _1766_ _1780_ _0907_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_108_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6306__A2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__A1 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7418_ _0241_ clknet_leaf_1_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _0172_ clknet_leaf_12_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3923__I _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5116__S _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6609__A3 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6490__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6174__C _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4556__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__A3 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7246__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3833__I _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5808__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7396__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6481__A1 _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3989__B _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__A4 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _0884_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6784__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6720_ _1990_ _2694_ _2044_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3932_ _3464_ _3465_ _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5709__B _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6651_ _2640_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3863_ _3213_ _3398_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6536__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ net53 _1632_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4547__A1 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6582_ as2650.stack\[7\]\[3\] _2579_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3794_ _3139_ as2650.r123\[0\]\[7\] _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4011__A3 _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5533_ _0837_ _1043_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _1497_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7203_ _0026_ clknet_leaf_58_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4415_ _0279_ _0608_ _0613_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5395_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7134_ _3083_ _3089_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4346_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7065_ _1428_ _1041_ _1015_ _1145_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4277_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6016_ _1984_ _2038_ _1575_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6472__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6224__B2 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6918_ _2896_ _2899_ _2705_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6849_ net35 _2832_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3918__I _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7269__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4002__A3 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6160__B1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3653__I as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5266__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__A1 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6463__B2 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4484__I _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__A2 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6766__A2 _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4529__A1 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__I _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4200_ as2650.holding_reg\[3\] _3560_ _0299_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4701__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5180_ _1296_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ _3579_ _3586_ _0268_ _3480_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_110_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6206__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6703_ _2676_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7411__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _3450_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4895_ _0401_ _0433_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__3738__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6509__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3991__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3846_ _3170_ _3172_ _3238_ _3241_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6634_ _0900_ _1299_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4062__C _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5193__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3777_ _3312_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6565_ _2498_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5732__A3 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3743__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4940__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5516_ _1048_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _3567_ _2464_ _2478_ _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__I _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5447_ _1504_ _0851_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5496__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5378_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4329_ _0463_ _0503_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7117_ _1675_ _0878_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__C _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7048_ _0605_ _3005_ _3010_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__A3 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3648__I _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3821__I3 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7173__A2 _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__I _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4479__I _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6436__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6987__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4998__A1 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4998__B2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3670__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3700_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3973__A2 _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4680_ _0820_ _0842_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _3149_ _3158_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6911__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _1411_ as2650.stack\[1\]\[11\] as2650.stack\[0\]\[11\] _0898_ _2364_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ _0944_ _1384_ _1388_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6281_ _2249_ _2297_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5232_ as2650.stack\[2\]\[11\] _1342_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5722__B _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4150__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5163_ as2650.stack\[3\]\[12\] _1290_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4114_ _3245_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5094_ _1250_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6978__A2 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ _3466_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6109__I _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5650__A2 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6553__B _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5938__B1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _2009_ _2011_ _2017_ _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _3510_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4878_ _1048_ _0447_ _3365_ _0815_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ _1579_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3829_ _3207_ _3364_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6548_ _1855_ _0549_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _1118_ _1854_ _2489_ _1204_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6666__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5469__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6418__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6969__A2 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7091__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4762__I _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3955__A2 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6910__C _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6354__B1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4904__A1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4937__I _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__A1 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7082__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4435__A3 _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A2 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4672__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5850_ _1873_ _1660_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4199__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A1 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1675_ _1812_ _1018_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3946__A2 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4732_ _3184_ _3188_ _3190_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7137__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3614_ as2650.cycle\[0\] _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6896__A1 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5699__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _1426_ _1893_ _2413_ _2414_ _1895_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4594_ _0535_ _0709_ _0752_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7382_ _0205_ clknet_leaf_58_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6333_ _2279_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4371__A2 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5008__I as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6264_ as2650.addr_buff\[0\] _1498_ _2278_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5215_ _1326_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6195_ as2650.pc\[6\] _1185_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3751__I _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5146_ _0955_ _1282_ _1284_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3882__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7073__A1 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5077_ _1216_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6820__A1 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4028_ _3561_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__I _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5979_ _3568_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3937__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4531__B _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5119__S _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6887__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4362__A2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6639__B2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6458__B _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__A2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5862__A2 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3873__A1 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7064__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6811__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3928__A2 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7119__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__I _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6878__A1 _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6212__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4353__A2 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__C _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5000_ as2650.overflow _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7055__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5605__A2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6951_ _2814_ _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _1013_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6882_ _2834_ _0599_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ _1854_ _1580_ _1858_ _1859_ _1571_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6030__A2 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3919__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ _1472_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4715_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4592__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5695_ _1731_ _0501_ _1704_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6869__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7434_ _0257_ clknet_leaf_18_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4646_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4577_ _0472_ _0727_ _0764_ _0710_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7365_ _0188_ clknet_leaf_38_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5961__I _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ as2650.pc\[10\] _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7296_ _0119_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6247_ _0857_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _1971_ _2196_ _2074_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7046__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__B _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ as2650.stack_ptr\[2\] _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5201__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A1 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6021__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__A1 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__A3 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__A4 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7128__I _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5532__A1 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4099__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3846__A1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4271__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6012__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6370__C _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__A2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__A1 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _0643_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5480_ _1535_ _1530_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4431_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7150_ _3072_ _3085_ _3102_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4362_ _0504_ _0519_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6101_ _0814_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6079__A2 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7081_ _0440_ _1701_ _3039_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4293_ _3383_ _0470_ _0496_ _3521_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _0832_ _2040_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _2333_ _2914_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _1760_ _2833_ _2224_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6003__A2 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1822_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6796_ _2739_ _2740_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5747_ _1761_ _1777_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5678_ _1620_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4317__A2 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7417_ _0240_ clknet_leaf_1_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5514__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5691__I _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7348_ _0171_ clknet_3_0_0_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _0102_ clknet_leaf_67_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__A4 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3828__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__B _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__CLK clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6490__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__I _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4005__A1 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5753__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6848__A4 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4859__A3 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__A2 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3819__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__B _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6481__A2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6365__C _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _0997_ _1062_ _1148_ _1150_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3931_ _3218_ _3428_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5992__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _3309_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _3187_ _3397_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ _1635_ _1644_ _1647_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6581_ _0944_ _2578_ _2582_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3793_ _3328_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_121_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5532_ _1452_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _1499_ _1501_ _1507_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _0025_ clknet_leaf_57_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4414_ as2650.r123\[1\]\[2\] _0610_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5394_ _0675_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7133_ _3326_ _3086_ _3088_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _0346_ _0530_ _0531_ _0389_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5016__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4276_ _0474_ _0475_ _0477_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7064_ _3326_ _3023_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4855__I _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _1987_ _1997_ _2036_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6472__A2 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6917_ _0980_ _2698_ _2898_ _2306_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6848_ net34 net51 net32 _2740_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5735__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _2635_ _2764_ _2765_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5127__S _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__B2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6185__C _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4226__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__I _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7213__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4529__A2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3844__I _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4130_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4061_ _0261_ _0264_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6454__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4465__A1 _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3807__A4 _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ net3 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6702_ net52 _2597_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4116__S _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3914_ _3134_ _3284_ _3449_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4894_ _0506_ _0558_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _2597_ _1425_ _1909_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3845_ _3324_ _3348_ _3379_ _3380_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5193__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _2510_ _0577_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6390__A1 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3776_ _3245_ _3311_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5515_ _1553_ _1561_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6495_ _0321_ _1554_ _2503_ _2504_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _3208_ _3194_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _3349_ _0863_ _0915_ _1428_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ _1570_ _1761_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4328_ _0458_ _0503_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4585__I _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ as2650.r123\[0\]\[7\] _3006_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4259_ _0357_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4456__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__S _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7236__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5956__A1 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7386__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__A1 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4695__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__A3 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6924__B _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4998__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3670__A2 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3973__A3 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3630_ _3159_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6372__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ as2650.stack\[1\]\[2\] _1385_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6280_ _0976_ _1886_ _2296_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ _0987_ _1341_ _1344_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__C _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _0991_ _1289_ _1293_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4113_ _0315_ _0316_ _3236_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5093_ as2650.stack\[5\]\[12\] _1249_ _1216_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4044_ _3314_ _3545_ _3577_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__I0 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6553__C _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5938__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3749__I _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ _0821_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _1113_ _1115_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4610__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _3304_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6616_ _2606_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3828_ _3173_ _3363_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5410__I0 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6547_ _1683_ _0535_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3759_ _3294_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_119_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _1413_ _3514_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6666__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5429_ _1175_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4429__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7091__A2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__C _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5929__A1 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A1 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6919__B _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6657__A2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7401__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3891__A2 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7082__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A3 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4840__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4800_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _1424_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _3398_ _0403_ _0914_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7137__A3 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__A2 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _2401_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6896__A2 _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3613_ _3148_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7381_ _0204_ clknet_3_2_0_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _0632_ _0778_ _0779_ _0664_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6332_ _2274_ _1528_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6263_ _2275_ _2279_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5214_ _1327_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6194_ as2650.pc\[7\] net2 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5320__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ as2650.stack\[3\]\[4\] _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3882__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _0976_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4863__I _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4027_ _3560_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4831__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _3328_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4929_ _3554_ _3493_ _3316_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_127_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5139__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__B _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__B _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5869__I _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__I0 _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7055__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4683__I _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _1538_ _2928_ _2929_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6802__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5901_ as2650.stack\[6\]\[0\] _1921_ _1922_ _1923_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6881_ _2861_ _2863_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5832_ _3306_ _1845_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6566__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5763_ _1737_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4041__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5694_ _1546_ _1714_ _1730_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7433_ _0256_ clknet_leaf_20_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4645_ _0672_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3963__S _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7364_ _0187_ clknet_leaf_54_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4576_ _0727_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6315_ _1240_ as2650.pc\[8\] _2251_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5463__B _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _0118_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6246_ _1902_ _2252_ _2262_ _1572_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6177_ _2072_ as2650.stack\[1\]\[6\] as2650.stack\[0\]\[6\] _1972_ _2196_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7046__A2 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5128_ _1271_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ as2650.pc\[4\] _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4280__A2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6309__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3791__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5532__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3672__I _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5296__A1 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6916__C _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7037__A2 _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5599__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4271__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3847__I _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5771__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3782__A1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _0621_ _3151_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4361_ _0558_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _2110_ _2118_ _2120_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _1700_ _0374_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4292_ _0364_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__A1 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ _0857_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5730__C _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _2334_ _2913_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4262__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _2609_ _2831_ _2847_ _1154_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6539__A1 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__B2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5815_ as2650.cycle\[5\] _1837_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6795_ _2770_ _2775_ _2780_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5211__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _1427_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5677_ _1712_ _1716_ _1717_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7416_ _0239_ clknet_leaf_2_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4628_ _0810_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6711__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5514__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__I0 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5193__B _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7347_ _0170_ clknet_leaf_11_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _0391_ _0687_ _0688_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7278_ _0101_ clknet_leaf_67_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _2210_ _2219_ _2246_ _2206_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6736__C _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7019__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6227__B1 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6950__A1 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5882__I _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6702__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4498__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__A4 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5269__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__B _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7292__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__I _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3930_ _3408_ _3433_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5992__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3861_ _3250_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5600_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ as2650.stack\[7\]\[2\] _2579_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5744__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6941__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3792_ _3137_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5462_ _1419_ _1514_ _1516_ _1081_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_7201_ _0024_ clknet_3_6_0_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4413_ _3530_ _0608_ _0612_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5393_ _1450_ _1459_ _1460_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7132_ _1720_ _3087_ _3080_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4344_ _3548_ _0532_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7063_ _3350_ _0637_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4275_ _3329_ as2650.r123_2\[1\]\[6\] _3338_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6556__C _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6014_ _1799_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _1241_ _2665_ _2897_ _2790_ _1939_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6291__C _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6847_ _2212_ _2830_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6778_ _2739_ _2674_ _2362_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5735__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3746__A1 _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5729_ _1761_ _0863_ _1762_ _1562_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__I _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6038__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4226__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5877__I _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A1 _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7176__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__B1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6923__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__I _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_51_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4162__A1 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7100__A1 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7100__B2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ _3587_ _0266_ _3430_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4217__A2 _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__I _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4962_ _1128_ _1129_ _1130_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _2681_ _2683_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3913_ net10 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3976__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7167__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ as2650.psl\[1\] _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3844_ _3320_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6914__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _2493_ _2566_ _2567_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3775_ _3304_ _3308_ _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_121_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7188__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ _1437_ _1008_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6494_ _1534_ _1123_ _1633_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5445_ _0810_ _1080_ _1000_ _0919_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_105_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4153__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _3214_ _0919_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7115_ _1125_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4327_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _0554_ _3005_ _3009_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4258_ _0397_ _0427_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4456__A2 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _3314_ _0362_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__A2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6220__I3 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6133__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4144__A1 _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4695__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4776__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7152__I _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__B1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5644__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6991__I _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3670__A3 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6940__B _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3855__I _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5230_ as2650.stack\[2\]\[10\] _1342_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4686__I _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ as2650.stack\[3\]\[11\] _1290_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3590__I _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4112_ _0317_ _3307_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ as2650.pc\[12\] _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5635__A1 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _3315_ _3553_ _3576_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__C _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__B _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5938__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _2012_ _2013_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6060__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _1114_ _3348_ _0464_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _1042_ _0843_ _0636_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3827_ _3174_ _3198_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6615_ _2605_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6546_ _1728_ _2455_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3758_ _3291_ _3293_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6115__A2 _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ _1129_ _1123_ _2486_ _2487_ _1412_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3689_ as2650.cycle\[3\] _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5428_ _0796_ _1478_ _1486_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5874__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ _3209_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4429__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _3284_ _0798_ _3449_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5929__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__B2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6760__B _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6354__A2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4117__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__A2 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4730_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _0844_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6345__A2 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6400_ _1249_ _2412_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3612_ _3135_ _3147_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7380_ _0203_ clknet_leaf_12_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4592_ _0549_ _0719_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6331_ _1707_ _2341_ _2343_ _2220_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _3280_ _2278_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7226__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5856__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5213_ _0951_ _1328_ _1333_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _2041_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5305__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _1274_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5608__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6805__B1 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7376__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _1236_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6281__A1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ _3556_ _3559_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6033__A1 _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5977_ _1955_ _1957_ _1999_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4595__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4928_ _0845_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _1023_ _1024_ _1027_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _2529_ _2530_ _2534_ _2535_ _2536_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_109_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__C _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5215__I _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3873__A3 as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6272__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6272__B2 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6811__A3 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__B1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__A2 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5834__B _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5689__I1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7399__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4510__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4964__I _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7055__A3 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6263__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _1921_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6880_ _2275_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6015__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5831_ _1708_ _1856_ _1857_ _1818_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_61_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__I _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6566__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4577__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5762_ _1776_ _1793_ _1794_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4713_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5693_ _1728_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7432_ _0255_ clknet_leaf_20_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4575_ _0758_ _0761_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7363_ _0186_ clknet_leaf_54_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6314_ _2249_ _2329_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7294_ _0117_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _2211_ _2261_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6176_ _1929_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5127_ as2650.stack\[4\]\[12\] _1249_ _1255_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5058_ _1223_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4265__B1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4009_ _3301_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6006__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A3 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6006__B2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4568__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4032__A3 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3791__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6493__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__A3 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6796__A2 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6548__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4559__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5220__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__A3 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3782__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__I _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _0449_ _0505_ _0507_ _0502_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ _0471_ _0314_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _0949_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__B _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4247__B1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _2300_ _2301_ _2855_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_81_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5739__B _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6863_ _2612_ _2833_ _2846_ _1742_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ _1515_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6794_ _2682_ _2778_ _2779_ _2617_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1765_ _1659_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5676_ _3580_ _1712_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7415_ _0238_ clknet_leaf_24_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4869__I _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4627_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6711__A2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__A1 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7346_ _0169_ clknet_leaf_11_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4558_ _0632_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4573__I1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7277_ _0100_ clknet_leaf_67_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4489_ _3216_ _0638_ _0674_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_89_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6475__A1 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _2217_ _2218_ _2236_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6159_ _2173_ _2177_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6227__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6227__B2 _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6778__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__I _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3948__I _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6702__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput40 net40 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5269__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6466__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__B _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6218__A1 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3860_ _3303_ _3314_ _3395_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ as2650.r0\[7\] _3145_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6941__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3755__A2 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ _0901_ _1517_ _1518_ _1014_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3593__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4412_ as2650.r123\[1\]\[1\] _0610_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7200_ _0023_ clknet_leaf_6_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5901__B1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ _0899_ _1449_ _0885_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7131_ _3084_ _0823_ _0805_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ _0536_ _0314_ _0364_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4180__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7062_ _0853_ _1099_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _3328_ as2650.r123\[1\]\[6\] _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _1995_ _2021_ _2032_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_98_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__A1 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5680__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6915_ _1760_ _2890_ _2310_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3768__I _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _2829_ _2817_ _2213_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6777_ _1226_ _2698_ _2763_ _1690_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5983__I _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3989_ _3416_ _3298_ _3523_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5735__A3 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ _1053_ _1056_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4599__I _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5659_ _1701_ _1636_ _1027_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_87_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4156__C1 _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7329_ _0152_ clknet_leaf_25_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A1 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6999__A2 _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3678__I _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5187__B2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__B1 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4162__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__A1 _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_20_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5133__I _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6673__B _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4972__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__A2 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3588__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4961_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _2684_ _2686_ _2688_ _1826_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3912_ _3396_ _3446_ _3447_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3976__A2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7167__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4892_ _3275_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5178__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6631_ _1439_ _0868_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3843_ _3169_ _3378_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4921__B _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__A2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3774_ _3309_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6562_ _1856_ _0600_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5513_ _1562_ _1018_ _1015_ _3261_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6493_ _1096_ _0741_ _2502_ _1158_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6678__A1 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5444_ _0655_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5350__A1 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4153__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _1436_ _1437_ _1438_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7114_ _3061_ _3070_ _3071_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4326_ _0517_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6139__I _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7045_ as2650.r123\[0\]\[6\] _3006_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4257_ _0357_ _0328_ _0371_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4456__A3 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4188_ _3521_ _0387_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7158__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6829_ _2659_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4916__A1 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4122__I _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4144__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6477__C _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5892__A2 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7094__B2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5644__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3655__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7101__C _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5837__B net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4907__A1 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__A1 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4967__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _0987_ _1289_ _1292_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4111_ as2650.cycle\[7\] _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7085__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5091_ _1248_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4042_ _3554_ _3322_ _3383_ _3575_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5635__A2 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5399__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5993_ _0818_ _2014_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6060__A2 _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _1114_ _0586_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4875_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6899__A1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6614_ _1631_ _2604_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6899__B2 _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3826_ _3361_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4374__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5571__A1 _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6545_ _1150_ _2538_ _2551_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3757_ as2650.ins_reg\[0\] _3292_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_88_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _0806_ _0726_ _3223_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3688_ _3153_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4877__I _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5427_ as2650.r123_2\[0\]\[7\] _1481_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4126__A2 _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3781__I _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ _1317_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4309_ _3478_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5289_ _0991_ _1376_ _1380_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4429__A3 _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7028_ _2997_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4062__A1 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5392__B _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4117__A2 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A2 _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7067__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6935__C _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7178__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__A3 _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4027__I _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6042__A2 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4660_ _0670_ _3272_ _0834_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3611_ _3141_ _3146_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4591_ _0536_ _0710_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _1243_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6261_ _2232_ _2276_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ as2650.stack\[2\]\[3\] _1329_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5856__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1234_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7058__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5143_ _1275_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5608__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6805__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ as2650.stack\[5\]\[7\] _1235_ _1227_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3619__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4025_ _3127_ _3557_ _3558_ _3130_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_65_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__B1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6033__A2 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _3505_ _1956_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7395__D _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ _3157_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5544__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3809_ _3344_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4347__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4789_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _0472_ _2463_ _1665_ _0381_ _2478_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_118_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _0806_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3858__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__A1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7320__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4283__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__B2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5406__I _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5838__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4274__A1 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5830_ _1742_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4026__A1 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ _1735_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5774__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3596__I _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5774__B2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4712_ as2650.stack_ptr\[1\] _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5692_ _0854_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7431_ _0254_ clknet_3_2_0_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ _0826_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4329__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _0185_ clknet_leaf_54_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4574_ _0481_ _0758_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5541__A4 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1241_ _1984_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7293_ _0116_ clknet_leaf_45_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7343__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5316__I _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6244_ _2259_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _1782_ _2187_ _2193_ _1779_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5126_ _1270_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ as2650.stack\[5\]\[3\] _1222_ _1217_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4265__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4265__B2 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5462__B1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4008_ _3523_ _3540_ _3541_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__S _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A4 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5765__A1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5959_ _0938_ _1936_ _1982_ _1695_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_71_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6190__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5226__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4130__I _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6766__B _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3846__A4 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6245__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4256__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5896__I _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4008__A1 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5756__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A1 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6181__B2 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4731__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ _3169_ _0472_ _0493_ _3321_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4247__A1 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6931_ _2814_ _2911_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _2840_ _2845_ _2769_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _1736_ _1841_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5747__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _1544_ _2682_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _3175_ _1309_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5675_ _1713_ _1714_ _1715_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7414_ _0237_ clknet_leaf_22_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6172__A1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _3183_ _3249_ _3190_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7345_ _0168_ clknet_leaf_11_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4557_ as2650.r0\[4\] _0690_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7276_ _0099_ clknet_leaf_67_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4488_ _0634_ _0680_ _0630_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6227_ _1429_ _2210_ _2244_ _1927_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6475__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4486__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6158_ _2085_ _2090_ _2133_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6227__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _1255_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4238__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6089_ _1974_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7239__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5738__A1 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__B1 _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7389__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput30 net30 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput41 net41 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6496__B _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4795__I _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__S0 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5729__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__B2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__I _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4401__A1 _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3790_ _3325_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3874__I _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__S _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6154__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5460_ _3212_ _1416_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _3448_ _0608_ _0611_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5391_ _1453_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7130_ _3084_ _3085_ _3077_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _3169_ _0374_ _0544_ _3321_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7061_ _1833_ _1578_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4273_ _3329_ as2650.r123_2\[0\]\[6\] _3333_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4468__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _2033_ _1987_ _2034_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
.ends

