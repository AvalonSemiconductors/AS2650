magic
tech gf180mcuD
magscale 1 5
timestamp 1701965447
<< obsm1 >>
rect 672 1538 74312 73569
<< metal2 >>
rect 1680 74600 1736 75000
rect 4144 74600 4200 75000
rect 6608 74600 6664 75000
rect 9072 74600 9128 75000
rect 11536 74600 11592 75000
rect 14000 74600 14056 75000
rect 16464 74600 16520 75000
rect 18928 74600 18984 75000
rect 21392 74600 21448 75000
rect 23856 74600 23912 75000
rect 26320 74600 26376 75000
rect 28784 74600 28840 75000
rect 31248 74600 31304 75000
rect 33712 74600 33768 75000
rect 36176 74600 36232 75000
rect 38640 74600 38696 75000
rect 41104 74600 41160 75000
rect 43568 74600 43624 75000
rect 46032 74600 46088 75000
rect 48496 74600 48552 75000
rect 50960 74600 51016 75000
rect 53424 74600 53480 75000
rect 55888 74600 55944 75000
rect 58352 74600 58408 75000
rect 60816 74600 60872 75000
rect 63280 74600 63336 75000
rect 65744 74600 65800 75000
rect 68208 74600 68264 75000
rect 70672 74600 70728 75000
rect 73136 74600 73192 75000
<< obsm2 >>
rect 630 74570 1650 74600
rect 1766 74570 4114 74600
rect 4230 74570 6578 74600
rect 6694 74570 9042 74600
rect 9158 74570 11506 74600
rect 11622 74570 13970 74600
rect 14086 74570 16434 74600
rect 16550 74570 18898 74600
rect 19014 74570 21362 74600
rect 21478 74570 23826 74600
rect 23942 74570 26290 74600
rect 26406 74570 28754 74600
rect 28870 74570 31218 74600
rect 31334 74570 33682 74600
rect 33798 74570 36146 74600
rect 36262 74570 38610 74600
rect 38726 74570 41074 74600
rect 41190 74570 43538 74600
rect 43654 74570 46002 74600
rect 46118 74570 48466 74600
rect 48582 74570 50930 74600
rect 51046 74570 53394 74600
rect 53510 74570 55858 74600
rect 55974 74570 58322 74600
rect 58438 74570 60786 74600
rect 60902 74570 63250 74600
rect 63366 74570 65714 74600
rect 65830 74570 68178 74600
rect 68294 74570 70642 74600
rect 70758 74570 73106 74600
rect 73222 74570 74186 74600
rect 630 1549 74186 74570
<< obsm3 >>
rect 625 1554 74191 73346
<< metal4 >>
rect 2224 1538 2384 73334
rect 9904 1538 10064 73334
rect 17584 1538 17744 73334
rect 25264 1538 25424 73334
rect 32944 1538 33104 73334
rect 40624 1538 40784 73334
rect 48304 1538 48464 73334
rect 55984 1538 56144 73334
rect 63664 1538 63824 73334
rect 71344 1538 71504 73334
<< obsm4 >>
rect 1806 2417 2194 73015
rect 2414 2417 9874 73015
rect 10094 2417 17554 73015
rect 17774 2417 25234 73015
rect 25454 2417 32914 73015
rect 33134 2417 40594 73015
rect 40814 2417 48274 73015
rect 48494 2417 55954 73015
rect 56174 2417 63634 73015
rect 63854 2417 71314 73015
rect 71534 2417 72170 73015
<< labels >>
rlabel metal2 s 1680 74600 1736 75000 6 DAC_clk
port 1 nsew signal output
rlabel metal2 s 6608 74600 6664 75000 6 DAC_dat_1
port 2 nsew signal output
rlabel metal2 s 9072 74600 9128 75000 6 DAC_dat_2
port 3 nsew signal output
rlabel metal2 s 4144 74600 4200 75000 6 DAC_le
port 4 nsew signal output
rlabel metal2 s 11536 74600 11592 75000 6 addr[0]
port 5 nsew signal input
rlabel metal2 s 14000 74600 14056 75000 6 addr[1]
port 6 nsew signal input
rlabel metal2 s 16464 74600 16520 75000 6 addr[2]
port 7 nsew signal input
rlabel metal2 s 18928 74600 18984 75000 6 addr[3]
port 8 nsew signal input
rlabel metal2 s 21392 74600 21448 75000 6 addr[4]
port 9 nsew signal input
rlabel metal2 s 23856 74600 23912 75000 6 addr[5]
port 10 nsew signal input
rlabel metal2 s 65744 74600 65800 75000 6 bus_cyc
port 11 nsew signal input
rlabel metal2 s 26320 74600 26376 75000 6 bus_in[0]
port 12 nsew signal input
rlabel metal2 s 28784 74600 28840 75000 6 bus_in[1]
port 13 nsew signal input
rlabel metal2 s 31248 74600 31304 75000 6 bus_in[2]
port 14 nsew signal input
rlabel metal2 s 33712 74600 33768 75000 6 bus_in[3]
port 15 nsew signal input
rlabel metal2 s 36176 74600 36232 75000 6 bus_in[4]
port 16 nsew signal input
rlabel metal2 s 38640 74600 38696 75000 6 bus_in[5]
port 17 nsew signal input
rlabel metal2 s 41104 74600 41160 75000 6 bus_in[6]
port 18 nsew signal input
rlabel metal2 s 43568 74600 43624 75000 6 bus_in[7]
port 19 nsew signal input
rlabel metal2 s 46032 74600 46088 75000 6 bus_out[0]
port 20 nsew signal output
rlabel metal2 s 48496 74600 48552 75000 6 bus_out[1]
port 21 nsew signal output
rlabel metal2 s 50960 74600 51016 75000 6 bus_out[2]
port 22 nsew signal output
rlabel metal2 s 53424 74600 53480 75000 6 bus_out[3]
port 23 nsew signal output
rlabel metal2 s 55888 74600 55944 75000 6 bus_out[4]
port 24 nsew signal output
rlabel metal2 s 58352 74600 58408 75000 6 bus_out[5]
port 25 nsew signal output
rlabel metal2 s 60816 74600 60872 75000 6 bus_out[6]
port 26 nsew signal output
rlabel metal2 s 63280 74600 63336 75000 6 bus_out[7]
port 27 nsew signal output
rlabel metal2 s 68208 74600 68264 75000 6 bus_we
port 28 nsew signal input
rlabel metal2 s 70672 74600 70728 75000 6 clk
port 29 nsew signal input
rlabel metal2 s 73136 74600 73192 75000 6 rst
port 30 nsew signal input
rlabel metal4 s 2224 1538 2384 73334 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 73334 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 73334 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 73334 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 73334 6 vdd
port 31 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 73334 6 vss
port 32 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 73334 6 vss
port 32 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 73334 6 vss
port 32 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 73334 6 vss
port 32 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 73334 6 vss
port 32 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 75000 75000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17197350
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/SID/runs/23_12_07_16_51/results/signoff/sid_top.magic.gds
string GDS_START 540520
<< end >>

