VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO boot_rom
  CLASS BLOCK ;
  FOREIGN boot_rom ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN WEb_raw
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 296.000 37.520 300.000 ;
    END
  END WEb_raw
  PIN bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 296.000 115.920 300.000 ;
    END
  END bus_in[0]
  PIN bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 296.000 127.120 300.000 ;
    END
  END bus_in[1]
  PIN bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 296.000 138.320 300.000 ;
    END
  END bus_in[2]
  PIN bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 296.000 149.520 300.000 ;
    END
  END bus_in[3]
  PIN bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 296.000 160.720 300.000 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 296.000 171.920 300.000 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 296.000 183.120 300.000 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 296.000 194.320 300.000 ;
    END
  END bus_in[7]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 296.000 205.520 300.000 ;
    END
  END bus_out[0]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 296.000 216.720 300.000 ;
    END
  END bus_out[1]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 296.000 227.920 300.000 ;
    END
  END bus_out[2]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 296.000 239.120 300.000 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 296.000 250.320 300.000 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 296.000 261.520 300.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 296.000 272.720 300.000 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 296.000 283.920 300.000 ;
    END
  END bus_out[7]
  PIN cs_port[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 81.760 296.000 82.320 300.000 ;
    END
  END cs_port[0]
  PIN cs_port[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 296.000 93.520 300.000 ;
    END
  END cs_port[1]
  PIN cs_port[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 296.000 104.720 300.000 ;
    END
  END cs_port[2]
  PIN le_hi_act
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 296.000 59.920 300.000 ;
    END
  END le_hi_act
  PIN le_lo_act
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 296.000 48.720 300.000 ;
    END
  END le_lo_act
  PIN ram_end[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.440 4.000 154.000 ;
    END
  END ram_end[0]
  PIN ram_end[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.040 4.000 243.600 ;
    END
  END ram_end[10]
  PIN ram_end[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END ram_end[11]
  PIN ram_end[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 4.000 261.520 ;
    END
  END ram_end[12]
  PIN ram_end[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.920 4.000 270.480 ;
    END
  END ram_end[13]
  PIN ram_end[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END ram_end[14]
  PIN ram_end[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 287.840 4.000 288.400 ;
    END
  END ram_end[15]
  PIN ram_end[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 4.000 162.960 ;
    END
  END ram_end[1]
  PIN ram_end[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END ram_end[2]
  PIN ram_end[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 4.000 180.880 ;
    END
  END ram_end[3]
  PIN ram_end[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END ram_end[4]
  PIN ram_end[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END ram_end[5]
  PIN ram_end[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END ram_end[6]
  PIN ram_end[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 4.000 216.720 ;
    END
  END ram_end[7]
  PIN ram_end[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 4.000 225.680 ;
    END
  END ram_end[8]
  PIN ram_end[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.080 4.000 234.640 ;
    END
  END ram_end[9]
  PIN ram_start[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.080 4.000 10.640 ;
    END
  END ram_start[0]
  PIN ram_start[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 4.000 100.240 ;
    END
  END ram_start[10]
  PIN ram_start[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 108.640 4.000 109.200 ;
    END
  END ram_start[11]
  PIN ram_start[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END ram_start[12]
  PIN ram_start[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 4.000 127.120 ;
    END
  END ram_start[13]
  PIN ram_start[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.520 4.000 136.080 ;
    END
  END ram_start[14]
  PIN ram_start[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END ram_start[15]
  PIN ram_start[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 4.000 19.600 ;
    END
  END ram_start[1]
  PIN ram_start[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 4.000 28.560 ;
    END
  END ram_start[2]
  PIN ram_start[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 4.000 37.520 ;
    END
  END ram_start[3]
  PIN ram_start[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 4.000 46.480 ;
    END
  END ram_start[4]
  PIN ram_start[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 4.000 55.440 ;
    END
  END ram_start[5]
  PIN ram_start[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 4.000 64.400 ;
    END
  END ram_start[6]
  PIN ram_start[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END ram_start[7]
  PIN ram_start[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 4.000 82.320 ;
    END
  END ram_start[8]
  PIN ram_start[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END ram_start[9]
  PIN rom_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 296.000 71.120 300.000 ;
    END
  END rom_enabled
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 296.000 26.320 300.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 296.000 15.120 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.210 ;
      LAYER Metal2 ;
        RECT 5.180 295.700 14.260 296.000 ;
        RECT 15.420 295.700 25.460 296.000 ;
        RECT 26.620 295.700 36.660 296.000 ;
        RECT 37.820 295.700 47.860 296.000 ;
        RECT 49.020 295.700 59.060 296.000 ;
        RECT 60.220 295.700 70.260 296.000 ;
        RECT 71.420 295.700 81.460 296.000 ;
        RECT 82.620 295.700 92.660 296.000 ;
        RECT 93.820 295.700 103.860 296.000 ;
        RECT 105.020 295.700 115.060 296.000 ;
        RECT 116.220 295.700 126.260 296.000 ;
        RECT 127.420 295.700 137.460 296.000 ;
        RECT 138.620 295.700 148.660 296.000 ;
        RECT 149.820 295.700 159.860 296.000 ;
        RECT 161.020 295.700 171.060 296.000 ;
        RECT 172.220 295.700 182.260 296.000 ;
        RECT 183.420 295.700 193.460 296.000 ;
        RECT 194.620 295.700 204.660 296.000 ;
        RECT 205.820 295.700 215.860 296.000 ;
        RECT 217.020 295.700 227.060 296.000 ;
        RECT 228.220 295.700 238.260 296.000 ;
        RECT 239.420 295.700 249.460 296.000 ;
        RECT 250.620 295.700 260.660 296.000 ;
        RECT 261.820 295.700 271.860 296.000 ;
        RECT 273.020 295.700 283.060 296.000 ;
        RECT 5.180 10.170 283.780 295.700 ;
      LAYER Metal3 ;
        RECT 4.300 287.540 280.470 288.260 ;
        RECT 4.000 279.740 280.470 287.540 ;
        RECT 4.300 278.580 280.470 279.740 ;
        RECT 4.000 270.780 280.470 278.580 ;
        RECT 4.300 269.620 280.470 270.780 ;
        RECT 4.000 261.820 280.470 269.620 ;
        RECT 4.300 260.660 280.470 261.820 ;
        RECT 4.000 252.860 280.470 260.660 ;
        RECT 4.300 251.700 280.470 252.860 ;
        RECT 4.000 243.900 280.470 251.700 ;
        RECT 4.300 242.740 280.470 243.900 ;
        RECT 4.000 234.940 280.470 242.740 ;
        RECT 4.300 233.780 280.470 234.940 ;
        RECT 4.000 225.980 280.470 233.780 ;
        RECT 4.300 224.820 280.470 225.980 ;
        RECT 4.000 217.020 280.470 224.820 ;
        RECT 4.300 215.860 280.470 217.020 ;
        RECT 4.000 208.060 280.470 215.860 ;
        RECT 4.300 206.900 280.470 208.060 ;
        RECT 4.000 199.100 280.470 206.900 ;
        RECT 4.300 197.940 280.470 199.100 ;
        RECT 4.000 190.140 280.470 197.940 ;
        RECT 4.300 188.980 280.470 190.140 ;
        RECT 4.000 181.180 280.470 188.980 ;
        RECT 4.300 180.020 280.470 181.180 ;
        RECT 4.000 172.220 280.470 180.020 ;
        RECT 4.300 171.060 280.470 172.220 ;
        RECT 4.000 163.260 280.470 171.060 ;
        RECT 4.300 162.100 280.470 163.260 ;
        RECT 4.000 154.300 280.470 162.100 ;
        RECT 4.300 153.140 280.470 154.300 ;
        RECT 4.000 145.340 280.470 153.140 ;
        RECT 4.300 144.180 280.470 145.340 ;
        RECT 4.000 136.380 280.470 144.180 ;
        RECT 4.300 135.220 280.470 136.380 ;
        RECT 4.000 127.420 280.470 135.220 ;
        RECT 4.300 126.260 280.470 127.420 ;
        RECT 4.000 118.460 280.470 126.260 ;
        RECT 4.300 117.300 280.470 118.460 ;
        RECT 4.000 109.500 280.470 117.300 ;
        RECT 4.300 108.340 280.470 109.500 ;
        RECT 4.000 100.540 280.470 108.340 ;
        RECT 4.300 99.380 280.470 100.540 ;
        RECT 4.000 91.580 280.470 99.380 ;
        RECT 4.300 90.420 280.470 91.580 ;
        RECT 4.000 82.620 280.470 90.420 ;
        RECT 4.300 81.460 280.470 82.620 ;
        RECT 4.000 73.660 280.470 81.460 ;
        RECT 4.300 72.500 280.470 73.660 ;
        RECT 4.000 64.700 280.470 72.500 ;
        RECT 4.300 63.540 280.470 64.700 ;
        RECT 4.000 55.740 280.470 63.540 ;
        RECT 4.300 54.580 280.470 55.740 ;
        RECT 4.000 46.780 280.470 54.580 ;
        RECT 4.300 45.620 280.470 46.780 ;
        RECT 4.000 37.820 280.470 45.620 ;
        RECT 4.300 36.660 280.470 37.820 ;
        RECT 4.000 28.860 280.470 36.660 ;
        RECT 4.300 27.700 280.470 28.860 ;
        RECT 4.000 19.900 280.470 27.700 ;
        RECT 4.300 18.740 280.470 19.900 ;
        RECT 4.000 10.940 280.470 18.740 ;
        RECT 4.300 10.220 280.470 10.940 ;
      LAYER Metal4 ;
        RECT 14.140 108.170 21.940 241.830 ;
        RECT 24.140 108.170 98.740 241.830 ;
        RECT 100.940 108.170 140.420 241.830 ;
  END
END boot_rom
END LIBRARY

