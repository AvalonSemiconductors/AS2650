// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire net90;
 wire clknet_leaf_0_wb_clk_i;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net91;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net92;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net93;
 wire net94;
 wire net79;
 wire net84;
 wire net80;
 wire net81;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net82;
 wire net83;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_2_1_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4261_ (.I(net26),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4262_ (.I(\as2650.ins_reg[0] ),
    .Z(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4263_ (.I(_3843_),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4264_ (.I(_3844_),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4265_ (.I(_3845_),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4266_ (.I(_3846_),
    .Z(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4267_ (.I(_3847_),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4268_ (.I(_3848_),
    .Z(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4269_ (.A1(\as2650.halted ),
    .A2(net10),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4270_ (.I(\as2650.psl[4] ),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4271_ (.I(_3851_),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4272_ (.I(_3852_),
    .Z(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4273_ (.I(_3853_),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4274_ (.I(_3854_),
    .Z(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4275_ (.I(_3855_),
    .Z(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4276_ (.I(\as2650.ins_reg[0] ),
    .Z(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4277_ (.I(\as2650.ins_reg[1] ),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4278_ (.A1(_3857_),
    .A2(_3858_),
    .ZN(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4279_ (.I(_3859_),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4280_ (.I(_3860_),
    .Z(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4281_ (.A1(_3856_),
    .A2(_3861_),
    .ZN(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4282_ (.A1(_3850_),
    .A2(_3862_),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4283_ (.I(_3863_),
    .Z(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4284_ (.I(_3864_),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4285_ (.I(\as2650.ins_reg[4] ),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4286_ (.I(_3866_),
    .Z(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4287_ (.I(\as2650.ins_reg[6] ),
    .Z(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4288_ (.I(_3868_),
    .ZN(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4289_ (.I(_3869_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4290_ (.A1(_3867_),
    .A2(_3870_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4291_ (.I(\as2650.ins_reg[3] ),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4292_ (.I(_3872_),
    .ZN(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4293_ (.I(_3873_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4294_ (.I(_3874_),
    .Z(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4295_ (.A1(\as2650.cycle[3] ),
    .A2(\as2650.cycle[2] ),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4296_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(\as2650.cycle[5] ),
    .A4(\as2650.cycle[4] ),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4297_ (.A1(_3876_),
    .A2(_3877_),
    .Z(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4298_ (.I(_3878_),
    .Z(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4299_ (.I(\as2650.cycle[1] ),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4300_ (.I(\as2650.cycle[0] ),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4301_ (.A1(_3880_),
    .A2(_3881_),
    .ZN(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4302_ (.A1(_3879_),
    .A2(_3882_),
    .ZN(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4303_ (.I(_3883_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4304_ (.A1(_3875_),
    .A2(_3884_),
    .ZN(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4305_ (.I(\as2650.ins_reg[4] ),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4306_ (.I(_3886_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4307_ (.I(_3887_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4308_ (.I(\as2650.cycle[7] ),
    .ZN(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4309_ (.I(\as2650.cycle[6] ),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4310_ (.I(\as2650.cycle[3] ),
    .ZN(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4311_ (.I(\as2650.cycle[2] ),
    .ZN(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4312_ (.A1(_3891_),
    .A2(_3892_),
    .ZN(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4313_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .A3(_3893_),
    .ZN(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4314_ (.I(\as2650.cycle[1] ),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4315_ (.I(\as2650.cycle[0] ),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4316_ (.A1(_3895_),
    .A2(_3896_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4317_ (.A1(_3890_),
    .A2(_3894_),
    .A3(_3897_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_3889_),
    .A2(_3898_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4319_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4320_ (.A1(_3888_),
    .A2(_3899_),
    .A3(_3900_),
    .ZN(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4321_ (.A1(_3871_),
    .A2(_3885_),
    .B(_3901_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4322_ (.I(_3874_),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4323_ (.I(_3876_),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4324_ (.I(_3877_),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4325_ (.A1(_3904_),
    .A2(_3905_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4326_ (.A1(\as2650.cycle[1] ),
    .A2(_3896_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4327_ (.A1(_3906_),
    .A2(_3907_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4328_ (.I(_3908_),
    .Z(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4329_ (.I(_3909_),
    .Z(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4330_ (.I(\as2650.ins_reg[2] ),
    .Z(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4331_ (.I(_3911_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4332_ (.I(\as2650.ins_reg[5] ),
    .Z(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4333_ (.I(_3913_),
    .Z(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4334_ (.I(\as2650.ins_reg[7] ),
    .Z(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4335_ (.I(_3915_),
    .ZN(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4336_ (.A1(_3868_),
    .A2(_3916_),
    .ZN(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4337_ (.A1(_3914_),
    .A2(_3917_),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4338_ (.A1(_3912_),
    .A2(_3887_),
    .A3(_3918_),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4339_ (.I(_3912_),
    .Z(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4340_ (.A1(\as2650.ins_reg[4] ),
    .A2(_3868_),
    .A3(\as2650.ins_reg[7] ),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4341_ (.A1(\as2650.ins_reg[5] ),
    .A2(_3921_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4342_ (.I(_3922_),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4343_ (.A1(_3920_),
    .A2(_3923_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4344_ (.A1(_3919_),
    .A2(_3924_),
    .ZN(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4345_ (.A1(_3903_),
    .A2(_3910_),
    .A3(_3925_),
    .ZN(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4346_ (.I(\as2650.addr_buff[7] ),
    .ZN(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4347_ (.I(_3889_),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4348_ (.I(_3894_),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4349_ (.A1(_3890_),
    .A2(_3929_),
    .A3(_3897_),
    .ZN(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4350_ (.A1(_3928_),
    .A2(_3930_),
    .ZN(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4351_ (.I(_3887_),
    .Z(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4352_ (.I(_3932_),
    .Z(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4353_ (.I(\as2650.addr_buff[5] ),
    .Z(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4354_ (.I(\as2650.addr_buff[6] ),
    .Z(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4355_ (.A1(_3934_),
    .A2(_3935_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4356_ (.A1(_3933_),
    .A2(_3936_),
    .ZN(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4357_ (.A1(_3927_),
    .A2(_3931_),
    .A3(_3937_),
    .ZN(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4358_ (.A1(_3902_),
    .A2(_3926_),
    .A3(_3938_),
    .ZN(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4359_ (.I(_3872_),
    .Z(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4360_ (.I(_3916_),
    .Z(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4361_ (.I(_3911_),
    .Z(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4362_ (.I(\as2650.ins_reg[4] ),
    .Z(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_3914_),
    .A2(_3943_),
    .ZN(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4364_ (.A1(_3942_),
    .A2(_3944_),
    .ZN(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4365_ (.A1(_3941_),
    .A2(_3945_),
    .ZN(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4366_ (.A1(\as2650.cycle[1] ),
    .A2(_3881_),
    .A3(_3878_),
    .ZN(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4367_ (.A1(_3940_),
    .A2(_3946_),
    .A3(_3947_),
    .ZN(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(_3864_),
    .A2(_3948_),
    .ZN(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4369_ (.I(_3949_),
    .Z(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4370_ (.I(_3856_),
    .Z(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4371_ (.I(_3951_),
    .Z(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4372_ (.I(\as2650.halted ),
    .Z(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4373_ (.I(_3953_),
    .ZN(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4374_ (.I(net10),
    .ZN(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4375_ (.A1(_3954_),
    .A2(_3955_),
    .ZN(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4376_ (.A1(_3952_),
    .A2(_3956_),
    .ZN(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4377_ (.I(_3896_),
    .Z(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4378_ (.I(\as2650.cycle[3] ),
    .Z(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4379_ (.A1(_3959_),
    .A2(_3892_),
    .ZN(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4380_ (.A1(_3905_),
    .A2(_3960_),
    .ZN(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4381_ (.A1(_3895_),
    .A2(_3961_),
    .ZN(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4382_ (.A1(_3958_),
    .A2(_3962_),
    .ZN(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4383_ (.A1(_3933_),
    .A2(_3963_),
    .ZN(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4384_ (.A1(\as2650.ins_reg[5] ),
    .A2(\as2650.ins_reg[6] ),
    .A3(\as2650.ins_reg[7] ),
    .ZN(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4385_ (.I(_3965_),
    .Z(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4386_ (.I(_3861_),
    .Z(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4387_ (.I(_3967_),
    .Z(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4388_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .ZN(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4389_ (.I(_3969_),
    .Z(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4390_ (.I(_3970_),
    .Z(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4391_ (.I(_3971_),
    .Z(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4392_ (.I(_3972_),
    .Z(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4393_ (.I(_3973_),
    .Z(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4394_ (.I(\as2650.idx_ctrl[1] ),
    .ZN(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4395_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4396_ (.A1(_3975_),
    .A2(_3976_),
    .ZN(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4397_ (.A1(_3968_),
    .A2(_3974_),
    .A3(_3977_),
    .ZN(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4398_ (.A1(_3957_),
    .A2(_3964_),
    .A3(_3966_),
    .A4(_3978_),
    .ZN(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4399_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4400_ (.I(_3980_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4401_ (.I(_3913_),
    .ZN(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4402_ (.I(\as2650.ins_reg[6] ),
    .Z(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4403_ (.A1(_3982_),
    .A2(_3983_),
    .A3(_3915_),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4404_ (.A1(_3943_),
    .A2(_3981_),
    .A3(_3984_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4405_ (.I(_3850_),
    .Z(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4406_ (.A1(_3986_),
    .A2(_3862_),
    .ZN(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4407_ (.A1(_3883_),
    .A2(_3987_),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4408_ (.A1(_3985_),
    .A2(_3988_),
    .ZN(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4409_ (.A1(_3950_),
    .A2(_3979_),
    .A3(_3989_),
    .ZN(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4410_ (.A1(_3865_),
    .A2(_3939_),
    .B(_3990_),
    .ZN(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4411_ (.A1(_3849_),
    .A2(_3991_),
    .Z(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4412_ (.I(_3979_),
    .Z(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4413_ (.I(_3913_),
    .Z(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4414_ (.I(_3994_),
    .Z(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4415_ (.A1(_3983_),
    .A2(_3915_),
    .ZN(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4416_ (.A1(_3995_),
    .A2(_3996_),
    .ZN(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4417_ (.I(_3997_),
    .Z(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4418_ (.I(\as2650.r0[0] ),
    .Z(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4419_ (.I(_3999_),
    .Z(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4420_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_3852_),
    .Z(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4421_ (.I(_4001_),
    .Z(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4422_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123_2[1][0] ),
    .S(_3852_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4423_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_3852_),
    .Z(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4424_ (.I0(_4000_),
    .I1(_4002_),
    .I2(_4003_),
    .I3(_4004_),
    .S0(_3843_),
    .S1(\as2650.ins_reg[1] ),
    .Z(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4425_ (.I(_4005_),
    .Z(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4426_ (.A1(\as2650.holding_reg[0] ),
    .A2(_3980_),
    .Z(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4427_ (.A1(_3969_),
    .A2(_4006_),
    .B(_4007_),
    .ZN(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4428_ (.I(\as2650.holding_reg[0] ),
    .Z(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4429_ (.I0(_4009_),
    .I1(_4006_),
    .S(_3980_),
    .Z(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4430_ (.A1(_4008_),
    .A2(_4010_),
    .Z(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4431_ (.I(_3915_),
    .Z(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4432_ (.A1(_3869_),
    .A2(_4012_),
    .ZN(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4433_ (.A1(_3982_),
    .A2(_4013_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4434_ (.I(_4014_),
    .Z(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4435_ (.I(\as2650.psl[3] ),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4436_ (.A1(_4016_),
    .A2(\as2650.carry ),
    .Z(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4437_ (.A1(_4017_),
    .A2(_4011_),
    .Z(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4438_ (.A1(_3983_),
    .A2(_3916_),
    .ZN(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4439_ (.I(_4019_),
    .Z(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4440_ (.I(_3982_),
    .Z(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(_4021_),
    .A2(_4020_),
    .ZN(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4442_ (.I(\as2650.carry ),
    .Z(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4443_ (.A1(\as2650.psl[3] ),
    .A2(_4023_),
    .ZN(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4444_ (.I(_4024_),
    .ZN(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4445_ (.A1(_4025_),
    .A2(_4011_),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4446_ (.I(_4010_),
    .Z(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4447_ (.A1(_3870_),
    .A2(_4012_),
    .ZN(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4448_ (.A1(_4021_),
    .A2(_4027_),
    .B(_4028_),
    .ZN(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4449_ (.A1(_4020_),
    .A2(_4008_),
    .B1(_4022_),
    .B2(_4026_),
    .C(_4029_),
    .ZN(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4450_ (.A1(_4015_),
    .A2(_4018_),
    .B(_4030_),
    .ZN(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4451_ (.I(_4005_),
    .Z(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4452_ (.A1(_4009_),
    .A2(_4032_),
    .ZN(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4453_ (.A1(_3918_),
    .A2(_4033_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4454_ (.A1(_3997_),
    .A2(_4034_),
    .ZN(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4455_ (.A1(_3998_),
    .A2(_4011_),
    .B1(_4031_),
    .B2(_4035_),
    .ZN(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4456_ (.I(_4036_),
    .Z(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4457_ (.A1(_3987_),
    .A2(_3938_),
    .ZN(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4458_ (.I(_4038_),
    .Z(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4459_ (.I(_4039_),
    .Z(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4460_ (.I(\as2650.addr_buff[6] ),
    .ZN(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4461_ (.A1(\as2650.addr_buff[5] ),
    .A2(_4041_),
    .ZN(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4462_ (.I(\as2650.addr_buff[5] ),
    .ZN(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4463_ (.A1(_4043_),
    .A2(_3935_),
    .ZN(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4464_ (.A1(_4042_),
    .A2(_4044_),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4465_ (.A1(_4032_),
    .A2(_4045_),
    .Z(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4466_ (.I(_4046_),
    .Z(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4467_ (.I(_3888_),
    .Z(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4468_ (.I(_3899_),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4469_ (.A1(_4048_),
    .A2(_4049_),
    .A3(_3900_),
    .ZN(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4470_ (.A1(_3864_),
    .A2(_4050_),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4471_ (.I(_4051_),
    .Z(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4472_ (.I(_4000_),
    .Z(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4473_ (.I(_4053_),
    .Z(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4474_ (.I(_4054_),
    .ZN(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4475_ (.A1(_3888_),
    .A2(_3984_),
    .ZN(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4476_ (.A1(_3974_),
    .A2(_4056_),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4477_ (.A1(_3909_),
    .A2(_3863_),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4478_ (.A1(_4057_),
    .A2(_4058_),
    .ZN(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4479_ (.I(_4059_),
    .Z(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4480_ (.I(_4060_),
    .Z(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4481_ (.I(_4059_),
    .Z(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4482_ (.I(net5),
    .Z(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4483_ (.I(_4063_),
    .Z(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4484_ (.I(_4064_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4485_ (.I(_3949_),
    .Z(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4486_ (.I(_4005_),
    .Z(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4487_ (.I(_4067_),
    .Z(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4488_ (.I(_4068_),
    .Z(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4489_ (.A1(_3921_),
    .A2(_4069_),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4490_ (.A1(_3950_),
    .A2(_4070_),
    .ZN(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4491_ (.A1(_3940_),
    .A2(_3919_),
    .ZN(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4492_ (.A1(_3988_),
    .A2(_4072_),
    .ZN(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4493_ (.I(_4073_),
    .Z(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4494_ (.A1(_4065_),
    .A2(_4066_),
    .B(_4071_),
    .C(_4074_),
    .ZN(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4495_ (.I(_3872_),
    .Z(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4496_ (.A1(_4076_),
    .A2(_3919_),
    .A3(_4058_),
    .ZN(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4497_ (.I(_4077_),
    .Z(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4498_ (.I(\as2650.r0[1] ),
    .Z(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4499_ (.I(_4079_),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4500_ (.I(_4080_),
    .ZN(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4501_ (.A1(_3844_),
    .A2(_3858_),
    .Z(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4502_ (.A1(_4081_),
    .A2(_4082_),
    .ZN(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4503_ (.A1(_3857_),
    .A2(_3858_),
    .Z(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4504_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_3854_),
    .Z(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4505_ (.A1(_4084_),
    .A2(_4085_),
    .Z(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4506_ (.A1(_3843_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4507_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(_3857_),
    .S1(_3854_),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4508_ (.A1(_4087_),
    .A2(_4088_),
    .Z(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4509_ (.A1(_4083_),
    .A2(_4086_),
    .A3(_4089_),
    .Z(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4510_ (.I(_4090_),
    .Z(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4511_ (.I(_4091_),
    .Z(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4512_ (.A1(_4076_),
    .A2(_3924_),
    .A3(_4058_),
    .ZN(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4513_ (.I(_4093_),
    .Z(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4514_ (.I(_4094_),
    .Z(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4515_ (.A1(_4078_),
    .A2(_4092_),
    .B(_4095_),
    .ZN(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4516_ (.I(\as2650.psl[3] ),
    .Z(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4517_ (.I(\as2650.r0[7] ),
    .Z(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_4098_),
    .Z(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4519_ (.A1(_4099_),
    .A2(_3861_),
    .ZN(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4520_ (.I(_4084_),
    .Z(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4521_ (.I(_4101_),
    .Z(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4522_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_3856_),
    .Z(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4523_ (.A1(_4102_),
    .A2(_4103_),
    .ZN(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4524_ (.I(_4087_),
    .Z(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4525_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_3845_),
    .S1(_3856_),
    .Z(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4526_ (.A1(_4105_),
    .A2(_4106_),
    .ZN(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4527_ (.A1(_4100_),
    .A2(_4104_),
    .A3(_4107_),
    .ZN(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4528_ (.I(_4108_),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4529_ (.I(_4109_),
    .Z(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4530_ (.A1(_4097_),
    .A2(_4110_),
    .B(_4017_),
    .ZN(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4531_ (.I(_4094_),
    .Z(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4532_ (.A1(_4075_),
    .A2(_4096_),
    .B1(_4111_),
    .B2(_4112_),
    .ZN(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4533_ (.A1(_4062_),
    .A2(_4113_),
    .ZN(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4534_ (.I(_4038_),
    .Z(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4535_ (.A1(_4055_),
    .A2(_4061_),
    .B(_4114_),
    .C(_4115_),
    .ZN(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4536_ (.A1(_4040_),
    .A2(_4047_),
    .B(_4052_),
    .C(_4116_),
    .ZN(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4537_ (.A1(_3865_),
    .A2(_4050_),
    .ZN(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4538_ (.I(_4118_),
    .Z(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4539_ (.A1(_3975_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4540_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_3976_),
    .ZN(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4541_ (.A1(_4120_),
    .A2(_4121_),
    .ZN(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4542_ (.A1(_4032_),
    .A2(_4122_),
    .Z(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4543_ (.I(_4123_),
    .Z(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4544_ (.A1(_4119_),
    .A2(_4124_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4545_ (.A1(_4117_),
    .A2(_4125_),
    .B(_3993_),
    .ZN(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4546_ (.A1(_3993_),
    .A2(_4037_),
    .B(_4126_),
    .ZN(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4547_ (.I(net10),
    .Z(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_3909_),
    .Z(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4549_ (.I(_4129_),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4550_ (.A1(_3957_),
    .A2(_4130_),
    .ZN(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4551_ (.A1(_3943_),
    .A2(_4019_),
    .ZN(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4552_ (.A1(_3994_),
    .A2(_4132_),
    .ZN(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4553_ (.A1(_3968_),
    .A2(_3973_),
    .A3(_4133_),
    .ZN(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4554_ (.I(_4134_),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4555_ (.A1(_4131_),
    .A2(_4135_),
    .ZN(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4556_ (.A1(_3964_),
    .A2(_3966_),
    .A3(_3978_),
    .ZN(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4557_ (.A1(_3952_),
    .A2(_3956_),
    .A3(_4137_),
    .ZN(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4558_ (.I(_3956_),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4559_ (.I(_3927_),
    .Z(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4560_ (.A1(_4140_),
    .A2(_3931_),
    .A3(_3937_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4561_ (.A1(_3902_),
    .A2(_3926_),
    .ZN(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4562_ (.A1(_4012_),
    .A2(_3944_),
    .ZN(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4563_ (.A1(_3911_),
    .A2(_3947_),
    .ZN(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4564_ (.A1(_3874_),
    .A2(_4143_),
    .A3(_4144_),
    .Z(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4565_ (.A1(_4141_),
    .A2(_4142_),
    .A3(_4145_),
    .B(_3862_),
    .ZN(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4566_ (.A1(_4139_),
    .A2(_4146_),
    .B(_3989_),
    .ZN(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4567_ (.A1(_4138_),
    .A2(_4147_),
    .ZN(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4568_ (.A1(_3848_),
    .A2(_4148_),
    .ZN(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4569_ (.A1(_4128_),
    .A2(_4136_),
    .A3(_4149_),
    .ZN(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4570_ (.I(_4150_),
    .Z(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4571_ (.A1(\as2650.r123[1][0] ),
    .A2(_4151_),
    .ZN(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4572_ (.I(_4054_),
    .Z(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4573_ (.I(_4136_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4574_ (.I(_4154_),
    .Z(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4575_ (.I(_4002_),
    .Z(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4576_ (.I(_4156_),
    .Z(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4577_ (.I(_4157_),
    .Z(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4578_ (.A1(_4153_),
    .A2(_4155_),
    .A3(_4158_),
    .ZN(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4579_ (.A1(_3992_),
    .A2(_4127_),
    .B(_4152_),
    .C(_4159_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_3992_),
    .Z(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_4138_),
    .Z(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4582_ (.I(_4161_),
    .Z(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4583_ (.I(_3994_),
    .Z(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4584_ (.I(_3996_),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4585_ (.A1(_4163_),
    .A2(_4164_),
    .Z(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4586_ (.A1(_4083_),
    .A2(_4086_),
    .A3(_4089_),
    .ZN(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4587_ (.A1(\as2650.holding_reg[1] ),
    .A2(_3970_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4588_ (.A1(_3970_),
    .A2(_4166_),
    .B(_4167_),
    .ZN(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4589_ (.A1(_4165_),
    .A2(_4168_),
    .ZN(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4590_ (.I(_3918_),
    .Z(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4591_ (.I(\as2650.holding_reg[1] ),
    .Z(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4592_ (.A1(_4171_),
    .A2(_4091_),
    .ZN(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4593_ (.A1(_4170_),
    .A2(_4172_),
    .ZN(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4594_ (.A1(\as2650.holding_reg[1] ),
    .A2(_4090_),
    .Z(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4595_ (.I(_4174_),
    .Z(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4596_ (.A1(_4008_),
    .A2(_4010_),
    .ZN(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4597_ (.A1(_4009_),
    .A2(_4068_),
    .B1(_4025_),
    .B2(_4176_),
    .ZN(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4598_ (.A1(_4175_),
    .A2(_4177_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4599_ (.A1(_4022_),
    .A2(_4178_),
    .ZN(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4600_ (.A1(_3995_),
    .A2(_4020_),
    .ZN(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4601_ (.A1(_4033_),
    .A2(_4027_),
    .B1(_4011_),
    .B2(_4017_),
    .ZN(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4602_ (.A1(_4175_),
    .A2(_4181_),
    .Z(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4603_ (.A1(_3995_),
    .A2(_4028_),
    .ZN(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4604_ (.I(_3981_),
    .Z(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4605_ (.I(_4166_),
    .Z(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4606_ (.A1(_4171_),
    .A2(_4184_),
    .ZN(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4607_ (.A1(_4184_),
    .A2(_4185_),
    .B(_4186_),
    .C(_4013_),
    .ZN(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4608_ (.A1(_4180_),
    .A2(_4182_),
    .B(_4183_),
    .C(_4187_),
    .ZN(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4609_ (.A1(_4171_),
    .A2(_4091_),
    .ZN(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4610_ (.A1(_4163_),
    .A2(_4189_),
    .ZN(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(_4028_),
    .A2(_4190_),
    .ZN(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4612_ (.A1(_4179_),
    .A2(_4188_),
    .B(_4191_),
    .ZN(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4613_ (.A1(_4173_),
    .A2(_4192_),
    .ZN(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4614_ (.A1(_4169_),
    .A2(_4193_),
    .Z(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4615_ (.I(_4194_),
    .Z(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4616_ (.I(_4080_),
    .Z(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4617_ (.I(_4196_),
    .Z(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4618_ (.I(_4197_),
    .Z(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4619_ (.I(_3989_),
    .Z(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4620_ (.A1(_3865_),
    .A2(_4141_),
    .ZN(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4621_ (.I(_4200_),
    .Z(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4622_ (.I(_4069_),
    .Z(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4623_ (.I(_4202_),
    .Z(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4624_ (.A1(_3913_),
    .A2(_3869_),
    .A3(_3916_),
    .ZN(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4625_ (.A1(_3886_),
    .A2(_4204_),
    .ZN(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4626_ (.A1(_3942_),
    .A2(_4205_),
    .ZN(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4627_ (.I(_4206_),
    .Z(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4628_ (.A1(_3903_),
    .A2(_4207_),
    .A3(_3988_),
    .ZN(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4629_ (.I(_4208_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4630_ (.I(_4073_),
    .Z(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4631_ (.I(_4210_),
    .Z(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4632_ (.I(\as2650.r0[2] ),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4633_ (.I(_4212_),
    .Z(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4634_ (.I(_4213_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4635_ (.A1(_4214_),
    .A2(_3859_),
    .ZN(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4636_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_3853_),
    .Z(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4637_ (.A1(_4084_),
    .A2(_4216_),
    .ZN(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4638_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_3843_),
    .S1(_3853_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4639_ (.A1(_4087_),
    .A2(_4218_),
    .ZN(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4640_ (.A1(_4215_),
    .A2(_4217_),
    .A3(_4219_),
    .ZN(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4641_ (.I(_4220_),
    .Z(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4642_ (.I(_4221_),
    .Z(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4643_ (.I(_4222_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4644_ (.I(net6),
    .ZN(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4645_ (.I(_4224_),
    .Z(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4646_ (.A1(_3864_),
    .A2(_4145_),
    .ZN(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(_4226_),
    .Z(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4648_ (.I(_4227_),
    .Z(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4649_ (.A1(\as2650.ins_reg[5] ),
    .A2(_3868_),
    .A3(\as2650.ins_reg[7] ),
    .Z(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4650_ (.A1(_3886_),
    .A2(_4229_),
    .ZN(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4651_ (.A1(_4068_),
    .A2(_4230_),
    .ZN(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4652_ (.A1(_3922_),
    .A2(_4068_),
    .Z(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4653_ (.A1(_4231_),
    .A2(_4232_),
    .ZN(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4654_ (.A1(_4185_),
    .A2(_4233_),
    .Z(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(_4227_),
    .A2(_4234_),
    .ZN(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4656_ (.A1(_4225_),
    .A2(_4228_),
    .B(_4235_),
    .C(_4074_),
    .ZN(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4657_ (.A1(_4211_),
    .A2(_4223_),
    .B(_4236_),
    .ZN(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4658_ (.A1(_4209_),
    .A2(_4237_),
    .ZN(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4659_ (.A1(_4203_),
    .A2(_4209_),
    .B(_4238_),
    .ZN(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4660_ (.A1(_4199_),
    .A2(_4239_),
    .ZN(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4661_ (.A1(_4198_),
    .A2(_4199_),
    .B(_4201_),
    .C(_4240_),
    .ZN(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4662_ (.A1(_3934_),
    .A2(_4041_),
    .ZN(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4663_ (.A1(_4067_),
    .A2(_4042_),
    .B(_4242_),
    .ZN(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4664_ (.A1(_4067_),
    .A2(_4166_),
    .A3(_4243_),
    .Z(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4665_ (.I(_4244_),
    .Z(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4666_ (.A1(_4040_),
    .A2(_4245_),
    .B(_4052_),
    .ZN(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4667_ (.A1(_3975_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4668_ (.A1(_4067_),
    .A2(_4120_),
    .B(_4247_),
    .ZN(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4669_ (.A1(_4202_),
    .A2(_4092_),
    .A3(_4248_),
    .Z(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4670_ (.I(_4138_),
    .Z(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4671_ (.A1(_4241_),
    .A2(_4246_),
    .B1(_4249_),
    .B2(_4052_),
    .C(_4250_),
    .ZN(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4672_ (.A1(_4162_),
    .A2(_4195_),
    .B(_4251_),
    .ZN(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4673_ (.I(_4150_),
    .Z(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4674_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_3851_),
    .Z(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4675_ (.I(_4254_),
    .Z(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4676_ (.I(_4255_),
    .Z(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4677_ (.I(_4256_),
    .Z(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4678_ (.A1(_4197_),
    .A2(_4053_),
    .A3(_4157_),
    .A4(_4257_),
    .ZN(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(_4257_),
    .Z(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4680_ (.I(_4259_),
    .Z(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4681_ (.A1(_4198_),
    .A2(_4158_),
    .B1(_4260_),
    .B2(_4153_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4682_ (.I(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4683_ (.A1(_4258_),
    .A2(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4684_ (.I(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4685_ (.A1(\as2650.r123[1][1] ),
    .A2(_4253_),
    .B1(_0287_),
    .B2(_4155_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4686_ (.A1(_4160_),
    .A2(_4252_),
    .B(_0288_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4687_ (.I(_4214_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4688_ (.I(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4689_ (.I(_4185_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4690_ (.I(\as2650.r0[3] ),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4691_ (.I(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4692_ (.I(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4693_ (.A1(_0294_),
    .A2(_3859_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4694_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_3854_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4695_ (.A1(_4101_),
    .A2(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4696_ (.I(_3853_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4697_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_3857_),
    .S1(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4698_ (.A1(_4105_),
    .A2(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4699_ (.A1(_0295_),
    .A2(_0297_),
    .A3(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4700_ (.I(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4701_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4702_ (.I(net7),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4703_ (.I(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4704_ (.I(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4705_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4706_ (.I(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4707_ (.A1(_4215_),
    .A2(_4217_),
    .A3(_4219_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4708_ (.I(_0309_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4709_ (.I(_0310_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4710_ (.I(_0311_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4711_ (.A1(_4005_),
    .A2(_4083_),
    .A3(_4086_),
    .A4(_4089_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4712_ (.I(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4713_ (.A1(_3866_),
    .A2(_3965_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4714_ (.I(_0315_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4715_ (.A1(_4092_),
    .A2(_4232_),
    .B1(_0314_),
    .B2(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4716_ (.A1(_0312_),
    .A2(_0317_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4717_ (.A1(_4227_),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4718_ (.A1(_0308_),
    .A2(_4228_),
    .B(_0319_),
    .C(_4210_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4719_ (.A1(_4211_),
    .A2(_0303_),
    .B(_0320_),
    .C(_4208_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4720_ (.A1(_0291_),
    .A2(_4209_),
    .B(_0321_),
    .C(_4199_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4721_ (.A1(_0290_),
    .A2(_4199_),
    .B(_4200_),
    .C(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4722_ (.A1(_4220_),
    .A2(_0313_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4723_ (.A1(_4044_),
    .A2(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4724_ (.I(_0309_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4725_ (.A1(_4083_),
    .A2(_4086_),
    .A3(_4089_),
    .B(_4006_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4726_ (.I(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4727_ (.A1(_0326_),
    .A2(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4728_ (.A1(_4045_),
    .A2(_4222_),
    .B1(_0329_),
    .B2(_4042_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4729_ (.A1(_0325_),
    .A2(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4730_ (.A1(_4040_),
    .A2(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4731_ (.A1(_4119_),
    .A2(_0323_),
    .A3(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4732_ (.I(_4051_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4733_ (.A1(_4121_),
    .A2(_0324_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4734_ (.A1(_4122_),
    .A2(_4222_),
    .B1(_0329_),
    .B2(_4120_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4735_ (.A1(_0335_),
    .A2(_0336_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4736_ (.A1(_0334_),
    .A2(_0337_),
    .B(_4161_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4737_ (.I(\as2650.holding_reg[2] ),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(_0339_),
    .A2(_4221_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4739_ (.A1(_0339_),
    .A2(_4221_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4740_ (.A1(_0340_),
    .A2(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4741_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4742_ (.A1(_4168_),
    .A2(_4172_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4743_ (.A1(_4174_),
    .A2(_4181_),
    .B(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4744_ (.A1(_0342_),
    .A2(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4745_ (.A1(_4189_),
    .A2(_4177_),
    .B(_4172_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4746_ (.A1(_0343_),
    .A2(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4747_ (.I(_4013_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4748_ (.A1(_4163_),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4749_ (.I(_4020_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4750_ (.A1(_0339_),
    .A2(_3980_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4751_ (.A1(_3981_),
    .A2(_0311_),
    .B(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4752_ (.I(_3917_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4753_ (.A1(_0351_),
    .A2(_0353_),
    .B(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4754_ (.A1(_4015_),
    .A2(_0346_),
    .B1(_0348_),
    .B2(_0350_),
    .C(_0355_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4755_ (.I(_4021_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4756_ (.I(_4028_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4757_ (.A1(_0358_),
    .A2(_0341_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4758_ (.A1(_0357_),
    .A2(_0340_),
    .B(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4759_ (.A1(_0356_),
    .A2(_0360_),
    .B(_3998_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4760_ (.A1(_3998_),
    .A2(_0343_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4761_ (.I(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4762_ (.A1(_0333_),
    .A2(_0338_),
    .B1(_0363_),
    .B2(_4162_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4763_ (.I(\as2650.psl[4] ),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4764_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(_0365_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4765_ (.I(_0366_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4766_ (.I(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4767_ (.I(_0368_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4768_ (.A1(_4053_),
    .A2(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4769_ (.A1(_0289_),
    .A2(_4157_),
    .B1(_4257_),
    .B2(_4196_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4770_ (.A1(_0289_),
    .A2(_4196_),
    .A3(_4156_),
    .A4(_4257_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4771_ (.A1(_0371_),
    .A2(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4772_ (.A1(_0370_),
    .A2(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4773_ (.A1(_4258_),
    .A2(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4774_ (.A1(\as2650.r123[1][2] ),
    .A2(_4253_),
    .B1(_0375_),
    .B2(_4154_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4775_ (.A1(_4160_),
    .A2(_0364_),
    .B(_0376_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4776_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_3976_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4777_ (.I(_4247_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4778_ (.A1(_0377_),
    .A2(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4779_ (.A1(_0295_),
    .A2(_0297_),
    .A3(_0300_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4780_ (.I(_0380_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4781_ (.I(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4782_ (.A1(_4032_),
    .A2(_4091_),
    .A3(_4221_),
    .A4(_0301_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4783_ (.A1(_0311_),
    .A2(_0328_),
    .B(_0381_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4784_ (.A1(_0383_),
    .A2(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4785_ (.A1(_0326_),
    .A2(_0313_),
    .A3(_0380_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4786_ (.A1(_0310_),
    .A2(_0314_),
    .B(_0381_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4787_ (.A1(_4121_),
    .A2(_0386_),
    .A3(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4788_ (.A1(_0379_),
    .A2(_0382_),
    .B1(_0385_),
    .B2(_0377_),
    .C(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4789_ (.I(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4790_ (.I(_0294_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4791_ (.I(_0312_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4792_ (.I(net8),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4793_ (.I(_0393_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4794_ (.I(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4795_ (.I(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4796_ (.I(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4797_ (.I(_0382_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4798_ (.A1(_0316_),
    .A2(_0311_),
    .A3(_0314_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4799_ (.A1(_4205_),
    .A2(_0312_),
    .A3(_0328_),
    .B(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4800_ (.A1(_0398_),
    .A2(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4801_ (.A1(_3950_),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4802_ (.A1(_0397_),
    .A2(_4066_),
    .B(_4074_),
    .C(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4803_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_3844_),
    .S1(_0298_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4804_ (.A1(_4105_),
    .A2(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4805_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_0298_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4806_ (.A1(_4101_),
    .A2(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4807_ (.I(\as2650.r0[4] ),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4808_ (.I(_0408_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4809_ (.I(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4810_ (.A1(_0410_),
    .A2(_3860_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4811_ (.A1(_0405_),
    .A2(_0407_),
    .A3(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4812_ (.I(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4813_ (.A1(_4078_),
    .A2(_0413_),
    .B(_4094_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4814_ (.A1(_4095_),
    .A2(_0392_),
    .B1(_0403_),
    .B2(_0414_),
    .C(_4060_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4815_ (.A1(_0391_),
    .A2(_4062_),
    .B(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4816_ (.A1(_4043_),
    .A2(_3935_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4817_ (.I(_4242_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4818_ (.A1(_0417_),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4819_ (.A1(_4044_),
    .A2(_0386_),
    .A3(_0387_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4820_ (.A1(_0419_),
    .A2(_0382_),
    .B1(_0385_),
    .B2(_0417_),
    .C(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4821_ (.I(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4822_ (.A1(_4039_),
    .A2(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4823_ (.A1(_4115_),
    .A2(_0416_),
    .B(_0423_),
    .C(_4118_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4824_ (.A1(_4119_),
    .A2(_0390_),
    .B(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4825_ (.I(_4165_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4826_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0302_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4827_ (.I(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4828_ (.I(\as2650.holding_reg[3] ),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4829_ (.A1(_0429_),
    .A2(_0302_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4830_ (.A1(_0428_),
    .A2(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4831_ (.I(_0431_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4832_ (.I(_4170_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4833_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3970_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4834_ (.A1(_3971_),
    .A2(_0310_),
    .B(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4835_ (.I(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4836_ (.A1(_0353_),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4837_ (.A1(_0342_),
    .A2(_0345_),
    .B(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4838_ (.A1(_0432_),
    .A2(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4839_ (.A1(_4189_),
    .A2(_4177_),
    .B(_0340_),
    .C(_4172_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4840_ (.A1(_0341_),
    .A2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4841_ (.A1(_0432_),
    .A2(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4842_ (.I(_3972_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4843_ (.I(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4844_ (.A1(_0444_),
    .A2(_0303_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4845_ (.I(_3981_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4846_ (.I(_0446_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4847_ (.A1(_0429_),
    .A2(_0447_),
    .B(_0351_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4848_ (.A1(_0350_),
    .A2(_0442_),
    .B1(_0445_),
    .B2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4849_ (.A1(_4180_),
    .A2(_0439_),
    .B(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4850_ (.A1(_0429_),
    .A2(_3971_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4851_ (.A1(_3971_),
    .A2(_0382_),
    .B(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4852_ (.A1(_0357_),
    .A2(_0452_),
    .B(_0358_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4853_ (.A1(_0433_),
    .A2(_0427_),
    .B1(_0450_),
    .B2(_0453_),
    .C(_0426_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4854_ (.A1(_0426_),
    .A2(_0432_),
    .B(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4855_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4856_ (.I0(_0425_),
    .I1(_0456_),
    .S(_4250_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4857_ (.I(_3909_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4858_ (.I(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4859_ (.I(_0459_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4860_ (.I(_3972_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4861_ (.A1(_3967_),
    .A2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4862_ (.A1(_3982_),
    .A2(_3887_),
    .A3(_4019_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4863_ (.A1(_0462_),
    .A2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4864_ (.A1(_3957_),
    .A2(_0460_),
    .A3(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4865_ (.I(_0465_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4866_ (.A1(_4258_),
    .A2(_0374_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4867_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(_0365_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4868_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4869_ (.A1(_4080_),
    .A2(_3999_),
    .A3(_0367_),
    .A4(_0469_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4870_ (.I(_0469_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4871_ (.I(_0471_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4872_ (.A1(_4196_),
    .A2(_0369_),
    .B1(_0472_),
    .B2(_4000_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4873_ (.A1(_0470_),
    .A2(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4874_ (.A1(_0294_),
    .A2(_4156_),
    .B1(_4256_),
    .B2(_0289_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4875_ (.A1(_0294_),
    .A2(_4214_),
    .A3(_4156_),
    .A4(_4256_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4876_ (.A1(_0475_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4877_ (.A1(_0474_),
    .A2(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4878_ (.I(_0372_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4879_ (.A1(_0370_),
    .A2(_0371_),
    .B(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4880_ (.A1(_0478_),
    .A2(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4881_ (.A1(_0467_),
    .A2(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4882_ (.A1(_0466_),
    .A2(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4883_ (.A1(\as2650.r123[1][3] ),
    .A2(_4151_),
    .B(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4884_ (.A1(_4160_),
    .A2(_0457_),
    .B(_0484_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4885_ (.I(\as2650.holding_reg[4] ),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4886_ (.A1(_0485_),
    .A2(_0461_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4887_ (.A1(_0446_),
    .A2(_0413_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4888_ (.A1(_0486_),
    .A2(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4889_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4890_ (.A1(_0426_),
    .A2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4891_ (.A1(_0485_),
    .A2(_0412_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4892_ (.A1(_4170_),
    .A2(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4893_ (.A1(_0405_),
    .A2(_0407_),
    .A3(_0411_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4894_ (.I(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4895_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4896_ (.A1(_0341_),
    .A2(_0440_),
    .B(_0428_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4897_ (.A1(_0430_),
    .A2(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4898_ (.A1(_0495_),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4899_ (.I(_0494_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4900_ (.A1(_0485_),
    .A2(_4184_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4901_ (.A1(_0447_),
    .A2(_0499_),
    .B(_0500_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4902_ (.A1(_0358_),
    .A2(_0489_),
    .B1(_0501_),
    .B2(_0349_),
    .C(_4170_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4903_ (.I(_0495_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_0427_),
    .A2(_0452_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4905_ (.A1(_0431_),
    .A2(_0438_),
    .B(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4906_ (.A1(_0503_),
    .A2(_0505_),
    .B(_4180_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4907_ (.A1(_0503_),
    .A2(_0505_),
    .B(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4908_ (.A1(_4022_),
    .A2(_0498_),
    .B(_0502_),
    .C(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4909_ (.A1(_0492_),
    .A2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4910_ (.A1(_0490_),
    .A2(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4911_ (.I(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4912_ (.I(_0417_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4913_ (.A1(_0310_),
    .A2(_0328_),
    .A3(_0381_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4914_ (.A1(_0494_),
    .A2(_0513_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4915_ (.A1(_0493_),
    .A2(_0386_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4916_ (.A1(_4045_),
    .A2(_0412_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4917_ (.A1(_0512_),
    .A2(_0514_),
    .B1(_0515_),
    .B2(_0418_),
    .C(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4918_ (.I(_0517_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4919_ (.I(_0410_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4920_ (.I(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4921_ (.I(_3858_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4922_ (.I(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4923_ (.A1(_3845_),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4924_ (.I0(\as2650.r123[1][5] ),
    .I1(\as2650.r123_2[1][5] ),
    .S(_3855_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4925_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123_2[0][5] ),
    .S(_0365_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4926_ (.I(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4927_ (.I(_0526_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4928_ (.I(_0527_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4929_ (.I(_3844_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4930_ (.A1(_0529_),
    .A2(_0521_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4931_ (.A1(_0523_),
    .A2(_0524_),
    .B1(_0528_),
    .B2(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4932_ (.I(\as2650.r0[5] ),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4933_ (.I(_0532_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4934_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_0298_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4935_ (.A1(_0533_),
    .A2(_3860_),
    .B1(_4101_),
    .B2(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4936_ (.A1(_0531_),
    .A2(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4937_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4938_ (.I(_0537_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4939_ (.I(_0538_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4940_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4941_ (.I(net9),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4942_ (.I(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4943_ (.I(_0542_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4944_ (.A1(_4222_),
    .A2(_0302_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4945_ (.A1(_0315_),
    .A2(_0314_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4946_ (.A1(_3923_),
    .A2(_0513_),
    .B1(_0544_),
    .B2(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4947_ (.A1(_0412_),
    .A2(_0546_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4948_ (.A1(_3949_),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4949_ (.A1(_0543_),
    .A2(_3950_),
    .B(_4210_),
    .C(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4950_ (.A1(_4074_),
    .A2(_0540_),
    .B(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4951_ (.A1(_4209_),
    .A2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4952_ (.A1(_4095_),
    .A2(_0303_),
    .B(_4060_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4953_ (.A1(_0520_),
    .A2(_4062_),
    .B1(_0551_),
    .B2(_0552_),
    .C(_4039_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4954_ (.A1(_4040_),
    .A2(_0518_),
    .B(_0553_),
    .C(_0334_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4955_ (.I(_0377_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4956_ (.A1(_0555_),
    .A2(_0514_),
    .B1(_0515_),
    .B2(_0378_),
    .C1(_0379_),
    .C2(_0499_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4957_ (.I(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4958_ (.A1(_4118_),
    .A2(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4959_ (.A1(_4161_),
    .A2(_0554_),
    .A3(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4960_ (.A1(_4162_),
    .A2(_0511_),
    .B(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4961_ (.I(\as2650.r0[1] ),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4962_ (.I(_0468_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4963_ (.A1(_0561_),
    .A2(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4964_ (.A1(_4213_),
    .A2(_0368_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4965_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123_2[0][4] ),
    .S(_0365_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4966_ (.I(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4967_ (.I(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4968_ (.I(_0567_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4969_ (.A1(_4000_),
    .A2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4970_ (.A1(_0563_),
    .A2(_0564_),
    .A3(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4971_ (.A1(_0293_),
    .A2(_4254_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4972_ (.A1(_0409_),
    .A2(_4001_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4973_ (.A1(_0470_),
    .A2(_0571_),
    .A3(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4974_ (.A1(_0570_),
    .A2(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4975_ (.A1(_0470_),
    .A2(_0473_),
    .A3(_0475_),
    .A4(_0476_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4976_ (.A1(_0476_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4977_ (.A1(_0574_),
    .A2(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4978_ (.A1(_0467_),
    .A2(_0481_),
    .A3(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4979_ (.A1(_0467_),
    .A2(_0481_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4980_ (.A1(_0478_),
    .A2(_0480_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4981_ (.A1(_0580_),
    .A2(_0577_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4982_ (.A1(_0579_),
    .A2(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4983_ (.A1(_0578_),
    .A2(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4984_ (.I(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4985_ (.A1(\as2650.r123[1][4] ),
    .A2(_4253_),
    .B1(_0584_),
    .B2(_4154_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4986_ (.A1(_4160_),
    .A2(_0560_),
    .B(_0585_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4987_ (.I(\as2650.holding_reg[5] ),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4988_ (.A1(_0586_),
    .A2(_0538_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4989_ (.A1(_0531_),
    .A2(_0535_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4990_ (.I(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4991_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4992_ (.A1(_0587_),
    .A2(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4993_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4994_ (.I(_0588_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4995_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4996_ (.I(_0447_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4997_ (.I(_0447_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4998_ (.A1(_0586_),
    .A2(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4999_ (.A1(_0595_),
    .A2(_0593_),
    .B(_0597_),
    .C(_0349_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5000_ (.A1(_0488_),
    .A2(_0491_),
    .B1(_0495_),
    .B2(_0505_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5001_ (.A1(_0592_),
    .A2(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5002_ (.A1(_0430_),
    .A2(_0495_),
    .A3(_0496_),
    .B(_0491_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5003_ (.A1(_0592_),
    .A2(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5004_ (.I(_4163_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5005_ (.A1(_0446_),
    .A2(_0538_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5006_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0446_),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5007_ (.A1(_0603_),
    .A2(_0605_),
    .B(_0354_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5008_ (.A1(_4015_),
    .A2(_0600_),
    .B1(_0602_),
    .B2(_0350_),
    .C(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5009_ (.A1(_0433_),
    .A2(_0594_),
    .B1(_0598_),
    .B2(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5010_ (.I(_3998_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5011_ (.I0(_0592_),
    .I1(_0608_),
    .S(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5012_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5013_ (.I(_0533_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5014_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5015_ (.I(_0499_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5016_ (.I(net1),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5017_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5018_ (.I(_0616_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5019_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5020_ (.A1(_0326_),
    .A2(_0327_),
    .A3(_0380_),
    .A4(_0493_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5021_ (.A1(_0326_),
    .A2(_0313_),
    .A3(_0380_),
    .A4(_0493_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5022_ (.A1(_3923_),
    .A2(_0619_),
    .B1(_0620_),
    .B2(_0316_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5023_ (.A1(_0593_),
    .A2(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5024_ (.A1(_4228_),
    .A2(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5025_ (.A1(_0618_),
    .A2(_4228_),
    .B(_0623_),
    .C(_4211_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5026_ (.I(\as2650.r0[6] ),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5027_ (.I(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5028_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5029_ (.A1(_0627_),
    .A2(_3860_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5030_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_3855_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5031_ (.A1(_4102_),
    .A2(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5032_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_3845_),
    .S1(_3855_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5033_ (.A1(_4105_),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5034_ (.A1(_0628_),
    .A2(_0630_),
    .A3(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5035_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5036_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5037_ (.A1(_4078_),
    .A2(_0635_),
    .B(_4095_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5038_ (.A1(_4112_),
    .A2(_0614_),
    .B1(_0624_),
    .B2(_0636_),
    .C(_4062_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5039_ (.A1(_0613_),
    .A2(_4061_),
    .B(_4115_),
    .C(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5040_ (.A1(_0537_),
    .A2(_0619_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5041_ (.A1(_0537_),
    .A2(_0620_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5042_ (.A1(_4045_),
    .A2(_0589_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5043_ (.A1(_0512_),
    .A2(_0639_),
    .B1(_0640_),
    .B2(_0418_),
    .C(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5044_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5045_ (.A1(_4201_),
    .A2(_0643_),
    .B(_4118_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5046_ (.A1(_4122_),
    .A2(_0589_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5047_ (.A1(_0555_),
    .A2(_0639_),
    .B1(_0640_),
    .B2(_0378_),
    .C(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5048_ (.A1(_0334_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5049_ (.A1(_0638_),
    .A2(_0644_),
    .B(_0647_),
    .C(_3993_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5050_ (.A1(_3993_),
    .A2(_0611_),
    .B(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5051_ (.A1(_0478_),
    .A2(_0480_),
    .A3(_0577_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5052_ (.A1(_0650_),
    .A2(_0578_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5053_ (.A1(_0574_),
    .A2(_0576_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5054_ (.A1(_0470_),
    .A2(_0571_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5055_ (.A1(_0653_),
    .A2(_0572_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5056_ (.A1(_0370_),
    .A2(_0563_),
    .A3(_0571_),
    .B(_0654_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5057_ (.A1(_0570_),
    .A2(_0573_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5058_ (.I(\as2650.r0[0] ),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5059_ (.A1(_0657_),
    .A2(_0527_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5060_ (.A1(_4079_),
    .A2(_0566_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5061_ (.A1(_0292_),
    .A2(_0367_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5062_ (.A1(_4213_),
    .A2(_0469_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5063_ (.A1(_0659_),
    .A2(_0660_),
    .A3(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5064_ (.A1(_0658_),
    .A2(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5065_ (.A1(_0532_),
    .A2(_4002_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5066_ (.A1(_0657_),
    .A2(_0471_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5067_ (.A1(_4080_),
    .A2(_0469_),
    .B1(_0567_),
    .B2(_0657_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5068_ (.A1(_0665_),
    .A2(_0659_),
    .B1(_0666_),
    .B2(_0564_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5069_ (.A1(_0409_),
    .A2(_4255_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5070_ (.A1(_0664_),
    .A2(_0667_),
    .A3(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5071_ (.A1(_0656_),
    .A2(_0663_),
    .A3(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5072_ (.A1(_0655_),
    .A2(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5073_ (.A1(_0652_),
    .A2(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5074_ (.A1(_0651_),
    .A2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5075_ (.A1(_0465_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5076_ (.A1(\as2650.r123[1][5] ),
    .A2(_4151_),
    .B(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5077_ (.A1(_3992_),
    .A2(_0649_),
    .B(_0675_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5078_ (.A1(_0628_),
    .A2(_0630_),
    .A3(_0632_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5079_ (.A1(\as2650.holding_reg[6] ),
    .A2(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5080_ (.I(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5081_ (.A1(_0587_),
    .A2(_0605_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5082_ (.A1(_0591_),
    .A2(_0599_),
    .B(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5083_ (.A1(_0678_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5084_ (.I(_0676_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5085_ (.I(\as2650.holding_reg[6] ),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5086_ (.A1(_0683_),
    .A2(_0443_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5087_ (.A1(_3974_),
    .A2(_0682_),
    .B(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5088_ (.A1(_0357_),
    .A2(_0685_),
    .B(_0358_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5089_ (.A1(_0586_),
    .A2(_0539_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5090_ (.A1(_0687_),
    .A2(_0601_),
    .B(_0587_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5091_ (.A1(_0677_),
    .A2(_0688_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5092_ (.I(_0682_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5093_ (.A1(_0683_),
    .A2(_0596_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5094_ (.A1(_0596_),
    .A2(_0690_),
    .B(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5095_ (.A1(_0350_),
    .A2(_0689_),
    .B1(_0692_),
    .B2(_0349_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5096_ (.A1(_4180_),
    .A2(_0681_),
    .B(_0686_),
    .C(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5097_ (.A1(_0683_),
    .A2(_0635_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5098_ (.A1(_0433_),
    .A2(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5099_ (.A1(_0609_),
    .A2(_0694_),
    .A3(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5100_ (.A1(_0609_),
    .A2(_0678_),
    .B(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5101_ (.A1(_0536_),
    .A2(_0620_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5102_ (.A1(_0676_),
    .A2(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5103_ (.A1(_0588_),
    .A2(_0619_),
    .A3(_0633_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5104_ (.A1(_0494_),
    .A2(_0383_),
    .A3(_0537_),
    .B(_0676_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5105_ (.A1(_0701_),
    .A2(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5106_ (.A1(_0555_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5107_ (.A1(_4122_),
    .A2(_0634_),
    .B1(_0700_),
    .B2(_4121_),
    .C(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5108_ (.I(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5109_ (.A1(_4044_),
    .A2(_0700_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5110_ (.A1(_0419_),
    .A2(_0682_),
    .B1(_0703_),
    .B2(_0512_),
    .C(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5111_ (.I(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5112_ (.I(_0627_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5113_ (.I(net2),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5114_ (.I(_0711_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5115_ (.I(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5116_ (.I(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5117_ (.A1(_0316_),
    .A2(_0538_),
    .A3(_0620_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5118_ (.A1(_3923_),
    .A2(_0589_),
    .A3(_0619_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5119_ (.A1(_0715_),
    .A2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5120_ (.A1(_0682_),
    .A2(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5121_ (.A1(_4226_),
    .A2(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5122_ (.A1(_0714_),
    .A2(_4227_),
    .B(_0719_),
    .C(_4210_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5123_ (.A1(_4077_),
    .A2(_4109_),
    .B(_4093_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5124_ (.A1(_4094_),
    .A2(_0539_),
    .B1(_0720_),
    .B2(_0721_),
    .C(_4059_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5125_ (.A1(_0710_),
    .A2(_4060_),
    .B(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5126_ (.A1(_4039_),
    .A2(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5127_ (.A1(_3865_),
    .A2(_3901_),
    .B1(_4115_),
    .B2(_0709_),
    .C(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5128_ (.A1(_0334_),
    .A2(_0706_),
    .B(_0725_),
    .C(_4161_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5129_ (.A1(_4250_),
    .A2(_0698_),
    .B(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5130_ (.A1(_0652_),
    .A2(_0671_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5131_ (.A1(_0651_),
    .A2(_0672_),
    .B(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5132_ (.I(_0670_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5133_ (.A1(_0663_),
    .A2(_0669_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5134_ (.A1(_0663_),
    .A2(_0669_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5135_ (.A1(_0656_),
    .A2(_0731_),
    .A3(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5136_ (.A1(_0655_),
    .A2(_0730_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5137_ (.A1(_0667_),
    .A2(_0668_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5138_ (.A1(_0667_),
    .A2(_0668_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5139_ (.A1(_0664_),
    .A2(_0735_),
    .A3(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5140_ (.A1(_0735_),
    .A2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5141_ (.A1(_0658_),
    .A2(_0662_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5142_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .S(_3851_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5143_ (.I(_0740_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5144_ (.A1(_3999_),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5145_ (.A1(_0561_),
    .A2(_0526_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5146_ (.I(_0740_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5147_ (.A1(_4079_),
    .A2(\as2650.r0[0] ),
    .A3(_0525_),
    .A4(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5148_ (.A1(_0742_),
    .A2(_0743_),
    .B(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(\as2650.r0[2] ),
    .A2(_0565_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5150_ (.A1(\as2650.r0[4] ),
    .A2(_0366_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5151_ (.A1(_0292_),
    .A2(_0562_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5152_ (.A1(_0747_),
    .A2(_0748_),
    .A3(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5153_ (.A1(_0746_),
    .A2(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5154_ (.A1(_4213_),
    .A2(_0562_),
    .B1(_0567_),
    .B2(_0561_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5155_ (.A1(_0563_),
    .A2(_0747_),
    .B1(_0752_),
    .B2(_0660_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5156_ (.A1(_0532_),
    .A2(_4255_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5157_ (.A1(_0625_),
    .A2(_4001_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5158_ (.A1(_0753_),
    .A2(_0754_),
    .A3(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5159_ (.A1(_0739_),
    .A2(_0751_),
    .A3(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5160_ (.A1(_0731_),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5161_ (.A1(_0738_),
    .A2(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5162_ (.A1(_0734_),
    .A2(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5163_ (.A1(_0729_),
    .A2(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5164_ (.A1(_0465_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5165_ (.A1(\as2650.r123[1][6] ),
    .A2(_4151_),
    .B(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5166_ (.A1(_3992_),
    .A2(_0727_),
    .B(_0763_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5167_ (.A1(_0734_),
    .A2(_0759_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5168_ (.A1(_0729_),
    .A2(_0760_),
    .B(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5169_ (.A1(_0738_),
    .A2(_0758_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5170_ (.A1(_0731_),
    .A2(_0757_),
    .B(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5171_ (.A1(_0612_),
    .A2(_4259_),
    .B(_0753_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5172_ (.A1(_0612_),
    .A2(_4259_),
    .A3(_0753_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5173_ (.A1(_0768_),
    .A2(_0755_),
    .B(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5174_ (.A1(_0739_),
    .A2(_0751_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5175_ (.A1(_0739_),
    .A2(_0751_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5176_ (.A1(_0771_),
    .A2(_0756_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5177_ (.A1(\as2650.r0[3] ),
    .A2(_0566_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5178_ (.A1(_0293_),
    .A2(_0471_),
    .B1(_0567_),
    .B2(_4214_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5179_ (.A1(_0661_),
    .A2(_0774_),
    .B1(_0775_),
    .B2(_0748_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5180_ (.A1(_0625_),
    .A2(_4255_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5181_ (.A1(_0776_),
    .A2(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5182_ (.A1(_4098_),
    .A2(_4002_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5183_ (.A1(_0778_),
    .A2(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5184_ (.A1(_0746_),
    .A2(_0750_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5185_ (.A1(\as2650.r0[5] ),
    .A2(_0367_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5186_ (.A1(_0408_),
    .A2(_0562_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5187_ (.A1(_0774_),
    .A2(_0782_),
    .A3(_0783_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5188_ (.A1(_4079_),
    .A2(_0744_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5189_ (.A1(_4212_),
    .A2(_0526_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5190_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_3851_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5191_ (.I(_0787_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5192_ (.A1(_0657_),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5193_ (.A1(_0785_),
    .A2(_0786_),
    .A3(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5194_ (.A1(_0745_),
    .A2(_0784_),
    .A3(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5195_ (.A1(_0781_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5196_ (.A1(_0780_),
    .A2(_0792_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5197_ (.A1(_0773_),
    .A2(_0793_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5198_ (.A1(_0770_),
    .A2(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5199_ (.A1(_0765_),
    .A2(_0767_),
    .A3(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5200_ (.A1(_4100_),
    .A2(_4104_),
    .A3(_4107_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5201_ (.A1(_4108_),
    .A2(_0701_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5202_ (.I(_0699_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5203_ (.A1(_0634_),
    .A2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5204_ (.A1(_0797_),
    .A2(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _5205_ (.A1(_0797_),
    .A2(_0419_),
    .B1(_0798_),
    .B2(_0512_),
    .C1(_0801_),
    .C2(_0418_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5206_ (.I(_0802_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5207_ (.I(_0635_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5208_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5209_ (.I(net3),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5210_ (.I(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5211_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5212_ (.A1(_4230_),
    .A2(_0634_),
    .A3(_0799_),
    .B1(_0701_),
    .B2(_4205_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5213_ (.A1(_4108_),
    .A2(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5214_ (.A1(_4066_),
    .A2(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5215_ (.A1(_0808_),
    .A2(_4066_),
    .B(_4211_),
    .C(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5216_ (.A1(\as2650.psl[3] ),
    .A2(_4069_),
    .B(_4017_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5217_ (.A1(_4078_),
    .A2(_0813_),
    .B(_4112_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5218_ (.A1(_4112_),
    .A2(_0805_),
    .B1(_0812_),
    .B2(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5219_ (.I(_4099_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5220_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5221_ (.A1(_0817_),
    .A2(_4061_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5222_ (.A1(_4061_),
    .A2(_0815_),
    .B(_0818_),
    .C(_4201_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5223_ (.A1(_4201_),
    .A2(_0803_),
    .B(_0819_),
    .C(_4119_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _5224_ (.A1(_0797_),
    .A2(_0379_),
    .B1(_0798_),
    .B2(_0555_),
    .C1(_0801_),
    .C2(_0378_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5225_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5226_ (.A1(_4052_),
    .A2(_0822_),
    .B(_4250_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5227_ (.I(\as2650.holding_reg[7] ),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5228_ (.I(_0797_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5229_ (.A1(_0824_),
    .A2(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5230_ (.A1(\as2650.holding_reg[7] ),
    .A2(_4109_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5231_ (.A1(_0826_),
    .A2(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5232_ (.I(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5233_ (.I(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5234_ (.A1(_0426_),
    .A2(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5235_ (.A1(_0678_),
    .A2(_0680_),
    .B1(_0685_),
    .B2(_0695_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5236_ (.A1(_0829_),
    .A2(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5237_ (.A1(_0677_),
    .A2(_0688_),
    .B(_0695_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5238_ (.A1(_0828_),
    .A2(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5239_ (.A1(_0824_),
    .A2(_0596_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5240_ (.A1(_0595_),
    .A2(_4109_),
    .B(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5241_ (.A1(_4022_),
    .A2(_0835_),
    .B1(_0837_),
    .B2(_0351_),
    .C(_4183_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5242_ (.A1(_4015_),
    .A2(_0833_),
    .B(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5243_ (.I(_0603_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5244_ (.A1(_0840_),
    .A2(_0826_),
    .B(_0354_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5245_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0433_),
    .A3(_4110_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5246_ (.A1(_0839_),
    .A2(_0841_),
    .B(_0842_),
    .C(_0609_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5247_ (.A1(_0831_),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5248_ (.A1(_0820_),
    .A2(_0823_),
    .B1(_0844_),
    .B2(_4162_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5249_ (.A1(\as2650.r123[1][7] ),
    .A2(_4253_),
    .B1(_0845_),
    .B2(_4149_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5250_ (.A1(_0466_),
    .A2(_0796_),
    .B(_0846_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5251_ (.I(_0521_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5252_ (.I(_0847_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5253_ (.I(_0848_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5254_ (.A1(_3886_),
    .A2(_3996_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5255_ (.A1(_3994_),
    .A2(_0462_),
    .A3(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5256_ (.A1(_3846_),
    .A2(_0522_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5257_ (.A1(_4184_),
    .A2(_0463_),
    .A3(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5258_ (.A1(_0851_),
    .A2(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5259_ (.I(_0854_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5260_ (.I(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5261_ (.A1(_4131_),
    .A2(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5262_ (.A1(_0848_),
    .A2(_4148_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5263_ (.A1(_4128_),
    .A2(_0857_),
    .A3(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5264_ (.I(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5265_ (.I(_0859_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5266_ (.A1(_3914_),
    .A2(_0850_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5267_ (.I(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5268_ (.A1(_3968_),
    .A2(_3974_),
    .A3(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5269_ (.I(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5270_ (.A1(_4131_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5271_ (.I(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5272_ (.A1(_4131_),
    .A2(_0856_),
    .B(_0465_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5273_ (.I(_0868_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5274_ (.I(_0851_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5275_ (.I(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5276_ (.I(\as2650.psu[0] ),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5277_ (.I(\as2650.psu[1] ),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5278_ (.I(_0873_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5279_ (.I(\as2650.psu[2] ),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5280_ (.A1(_0872_),
    .A2(_0874_),
    .B(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5281_ (.A1(_0872_),
    .A2(_0873_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5282_ (.A1(\as2650.psu[2] ),
    .A2(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5283_ (.A1(_0876_),
    .A2(_0878_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5284_ (.I(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5285_ (.I(_0880_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5286_ (.I(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5287_ (.I(\as2650.psu[0] ),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5288_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5289_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5290_ (.I(\as2650.psu[1] ),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5291_ (.I(_0886_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5292_ (.I0(\as2650.stack[7][8] ),
    .I1(\as2650.stack[4][8] ),
    .I2(\as2650.stack[5][8] ),
    .I3(\as2650.stack[6][8] ),
    .S0(_0885_),
    .S1(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5293_ (.A1(\as2650.psu[0] ),
    .A2(_0886_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5294_ (.I(_0877_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5295_ (.A1(_0889_),
    .A2(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5296_ (.I(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5297_ (.I(_0892_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5298_ (.I(_0893_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5299_ (.I(_0874_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5300_ (.I(_0895_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5301_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5302_ (.I(_0872_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5303_ (.I(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5304_ (.I(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5305_ (.I(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5306_ (.A1(_0897_),
    .A2(\as2650.stack[1][8] ),
    .B1(\as2650.stack[0][8] ),
    .B2(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5307_ (.I(_0875_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5308_ (.I(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5309_ (.I(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5310_ (.I(_0889_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5311_ (.I(_0906_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5313_ (.A1(_0905_),
    .A2(\as2650.stack[3][8] ),
    .B1(\as2650.stack[2][8] ),
    .B2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5314_ (.I(_0881_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5315_ (.A1(_0894_),
    .A2(_0902_),
    .B(_0909_),
    .C(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5316_ (.A1(_0882_),
    .A2(_0888_),
    .B(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5317_ (.A1(_0871_),
    .A2(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5318_ (.A1(_4153_),
    .A2(_0867_),
    .B(_0869_),
    .C(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5319_ (.A1(_0861_),
    .A2(_0914_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5320_ (.A1(\as2650.r123[0][0] ),
    .A2(_0860_),
    .B(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5321_ (.A1(_0849_),
    .A2(_3991_),
    .A3(_4127_),
    .B(_0916_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5322_ (.I(_0866_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5323_ (.I(_0881_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5324_ (.I0(\as2650.stack[7][9] ),
    .I1(\as2650.stack[4][9] ),
    .I2(\as2650.stack[5][9] ),
    .I3(\as2650.stack[6][9] ),
    .S0(_0885_),
    .S1(_0887_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5325_ (.I(_0907_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5326_ (.I(_0896_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5327_ (.A1(_0921_),
    .A2(\as2650.stack[1][9] ),
    .B1(\as2650.stack[0][9] ),
    .B2(_0901_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5328_ (.A1(_0920_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5329_ (.I(_0904_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5330_ (.A1(_0924_),
    .A2(\as2650.stack[3][9] ),
    .B1(\as2650.stack[2][9] ),
    .B2(_0908_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5331_ (.A1(_0918_),
    .A2(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5332_ (.A1(_0918_),
    .A2(_0919_),
    .B1(_0923_),
    .B2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5333_ (.A1(_0871_),
    .A2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5334_ (.A1(_4198_),
    .A2(_0917_),
    .B(_0868_),
    .C(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5335_ (.A1(_0859_),
    .A2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5336_ (.A1(\as2650.r123[0][1] ),
    .A2(_0860_),
    .B(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5337_ (.A1(_0849_),
    .A2(_3991_),
    .A3(_4252_),
    .B(_0931_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5338_ (.I(\as2650.r123[0][2] ),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5339_ (.I(_0859_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5340_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5341_ (.I(_0364_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5342_ (.I(_0858_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5343_ (.I(_0910_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5344_ (.I(_0885_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5345_ (.I(_0886_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5346_ (.I0(\as2650.stack[7][10] ),
    .I1(\as2650.stack[4][10] ),
    .I2(\as2650.stack[5][10] ),
    .I3(\as2650.stack[6][10] ),
    .S0(_0938_),
    .S1(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5347_ (.I(_0907_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5348_ (.I(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5349_ (.I(_0900_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5350_ (.A1(_0921_),
    .A2(\as2650.stack[1][10] ),
    .B1(\as2650.stack[0][10] ),
    .B2(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(_0942_),
    .A2(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5352_ (.A1(_0924_),
    .A2(\as2650.stack[3][10] ),
    .B1(\as2650.stack[2][10] ),
    .B2(_0920_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5353_ (.A1(_0882_),
    .A2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5354_ (.A1(_0937_),
    .A2(_0940_),
    .B1(_0945_),
    .B2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5355_ (.I(_0290_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5356_ (.A1(_0949_),
    .A2(_0866_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5357_ (.A1(_4136_),
    .A2(_0857_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5358_ (.A1(_0871_),
    .A2(_0948_),
    .B(_0950_),
    .C(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5359_ (.A1(_0935_),
    .A2(_0936_),
    .B(_0933_),
    .C(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5360_ (.A1(_0932_),
    .A2(_0934_),
    .B(_0953_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5361_ (.I(\as2650.r123[0][3] ),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5362_ (.I(_0457_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5363_ (.I0(\as2650.stack[7][11] ),
    .I1(\as2650.stack[4][11] ),
    .I2(\as2650.stack[5][11] ),
    .I3(\as2650.stack[6][11] ),
    .S0(_0884_),
    .S1(_0887_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5364_ (.A1(_0897_),
    .A2(\as2650.stack[1][11] ),
    .B1(\as2650.stack[0][11] ),
    .B2(_0901_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5365_ (.A1(_0941_),
    .A2(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5366_ (.A1(_0905_),
    .A2(\as2650.stack[3][11] ),
    .B1(\as2650.stack[2][11] ),
    .B2(_0908_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5367_ (.A1(_0910_),
    .A2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5368_ (.A1(_0918_),
    .A2(_0956_),
    .B1(_0958_),
    .B2(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5369_ (.I(_0391_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5370_ (.A1(_0962_),
    .A2(_0917_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5371_ (.A1(_0867_),
    .A2(_0961_),
    .B(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5372_ (.A1(_0955_),
    .A2(_0936_),
    .B1(_0869_),
    .B2(_0964_),
    .C(_0861_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5373_ (.A1(_0954_),
    .A2(_0934_),
    .B(_0965_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5374_ (.I(\as2650.r123[0][4] ),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5375_ (.I(_0870_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5376_ (.I0(\as2650.stack[7][12] ),
    .I1(\as2650.stack[4][12] ),
    .I2(\as2650.stack[5][12] ),
    .I3(\as2650.stack[6][12] ),
    .S0(_0938_),
    .S1(_0939_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5377_ (.A1(_0921_),
    .A2(\as2650.stack[1][12] ),
    .B1(\as2650.stack[0][12] ),
    .B2(_0943_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5378_ (.A1(_0942_),
    .A2(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5379_ (.A1(_0924_),
    .A2(\as2650.stack[3][12] ),
    .B1(\as2650.stack[2][12] ),
    .B2(_0920_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5380_ (.A1(_0882_),
    .A2(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5381_ (.A1(_0937_),
    .A2(_0968_),
    .B1(_0970_),
    .B2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5382_ (.A1(_0519_),
    .A2(_0917_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5383_ (.A1(_0967_),
    .A2(_0973_),
    .B(_0974_),
    .C(_0951_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5384_ (.A1(_0933_),
    .A2(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5385_ (.A1(_0849_),
    .A2(_4148_),
    .A3(_0560_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5386_ (.A1(_0966_),
    .A2(_0860_),
    .B1(_0976_),
    .B2(_0977_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5387_ (.I(\as2650.r123[0][5] ),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5388_ (.I(_0649_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5389_ (.I0(\as2650.stack[7][13] ),
    .I1(\as2650.stack[4][13] ),
    .I2(\as2650.stack[5][13] ),
    .I3(\as2650.stack[6][13] ),
    .S0(_0884_),
    .S1(_0886_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5390_ (.A1(_0897_),
    .A2(\as2650.stack[1][13] ),
    .B1(\as2650.stack[0][13] ),
    .B2(_0901_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5391_ (.A1(_0941_),
    .A2(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5392_ (.A1(_0905_),
    .A2(\as2650.stack[3][13] ),
    .B1(\as2650.stack[2][13] ),
    .B2(_0908_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5393_ (.A1(_0910_),
    .A2(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5394_ (.A1(_0918_),
    .A2(_0980_),
    .B1(_0982_),
    .B2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5395_ (.I(_0613_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5396_ (.A1(_0986_),
    .A2(_0917_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5397_ (.A1(_0867_),
    .A2(_0985_),
    .B(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5398_ (.A1(_0979_),
    .A2(_0936_),
    .B1(_0869_),
    .B2(_0988_),
    .C(_0861_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5399_ (.A1(_0978_),
    .A2(_0934_),
    .B(_0989_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5400_ (.I(\as2650.r123[0][6] ),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5401_ (.I(_0727_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5402_ (.I0(\as2650.stack[7][14] ),
    .I1(\as2650.stack[4][14] ),
    .I2(\as2650.stack[5][14] ),
    .I3(\as2650.stack[6][14] ),
    .S0(_0938_),
    .S1(_0939_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5403_ (.A1(_0921_),
    .A2(\as2650.stack[1][14] ),
    .B1(\as2650.stack[0][14] ),
    .B2(_0943_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5404_ (.A1(_0920_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5405_ (.A1(_0924_),
    .A2(\as2650.stack[3][14] ),
    .B1(\as2650.stack[2][14] ),
    .B2(_0941_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5406_ (.A1(_0882_),
    .A2(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5407_ (.A1(_0937_),
    .A2(_0992_),
    .B1(_0994_),
    .B2(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5408_ (.I(_0710_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5409_ (.A1(_0998_),
    .A2(_0866_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5410_ (.A1(_0867_),
    .A2(_0997_),
    .B(_0999_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5411_ (.A1(_0991_),
    .A2(_0858_),
    .B1(_0869_),
    .B2(_1000_),
    .C(_0861_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5412_ (.A1(_0990_),
    .A2(_0934_),
    .B(_1001_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5413_ (.I(\as2650.r123[0][7] ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5414_ (.I(_0817_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5415_ (.I(_1003_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5416_ (.A1(_1004_),
    .A2(_0967_),
    .A3(_0951_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5417_ (.A1(_0845_),
    .A2(_0936_),
    .B(_0933_),
    .C(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5418_ (.A1(_1002_),
    .A2(_0860_),
    .B(_1006_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5419_ (.I(_3883_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5420_ (.A1(_3973_),
    .A2(_0530_),
    .A3(_0862_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5421_ (.A1(_3956_),
    .A2(_1007_),
    .A3(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5422_ (.I(_1009_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5423_ (.A1(_0900_),
    .A2(_1010_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5424_ (.I(_1009_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5425_ (.I(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5426_ (.I(_0889_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5427_ (.A1(_1014_),
    .A2(_0890_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5428_ (.A1(_1015_),
    .A2(_1010_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5429_ (.A1(_0897_),
    .A2(_1013_),
    .B(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5430_ (.I(\as2650.psu[2] ),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5431_ (.I(_0876_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5432_ (.A1(_1019_),
    .A2(_0878_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5433_ (.I(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5434_ (.A1(_1021_),
    .A2(_1012_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5435_ (.A1(_1018_),
    .A2(_1012_),
    .B(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5436_ (.I(_3920_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5437_ (.I(_3906_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5438_ (.I(_3895_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5439_ (.I(_3881_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5440_ (.A1(_1026_),
    .A2(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5441_ (.A1(_1025_),
    .A2(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5442_ (.A1(_1024_),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5443_ (.I(_3880_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5444_ (.I(_3905_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5445_ (.A1(_1031_),
    .A2(_1032_),
    .A3(_3960_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5446_ (.A1(_1027_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5447_ (.A1(\as2650.addr_buff[7] ),
    .A2(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5448_ (.I(_3963_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5449_ (.I(_3892_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5450_ (.A1(_3959_),
    .A2(_1037_),
    .A3(_3880_),
    .A4(_3905_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5451_ (.I(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5452_ (.A1(_1027_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(_1036_),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5454_ (.A1(_1035_),
    .A2(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5455_ (.I(_3940_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5456_ (.A1(_3873_),
    .A2(_3867_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5457_ (.A1(_4019_),
    .A2(_4102_),
    .A3(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5458_ (.I(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5459_ (.A1(_1043_),
    .A2(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5460_ (.I(_3888_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5461_ (.A1(_1048_),
    .A2(_4014_),
    .B(_4143_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5462_ (.A1(_1030_),
    .A2(_1042_),
    .B(_1047_),
    .C(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5463_ (.I(_3963_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5464_ (.I(_3942_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5465_ (.A1(_3846_),
    .A2(_0521_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5466_ (.A1(_3872_),
    .A2(_3943_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5467_ (.A1(_4013_),
    .A2(_1053_),
    .A3(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5468_ (.A1(_1052_),
    .A2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5469_ (.I(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5470_ (.I(_1008_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5471_ (.I(_3884_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5472_ (.A1(_0357_),
    .A2(_1051_),
    .A3(_1057_),
    .B1(_1058_),
    .B2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5473_ (.A1(_1050_),
    .A2(_1060_),
    .B(_3986_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5474_ (.I(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5475_ (.A1(_1023_),
    .A2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5476_ (.A1(_1017_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5477_ (.A1(_1011_),
    .A2(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5478_ (.I(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5479_ (.I(_1066_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5480_ (.I(\as2650.pc[0] ),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5481_ (.I(_1068_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5482_ (.I(_1069_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5483_ (.I(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5484_ (.I(_4055_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5485_ (.I(_1013_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5486_ (.I(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5487_ (.I0(_1071_),
    .I1(_1072_),
    .S(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5488_ (.I(_1075_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5489_ (.I(_1065_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5490_ (.I(_1077_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5491_ (.A1(\as2650.stack[0][0] ),
    .A2(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5492_ (.A1(_1067_),
    .A2(_1076_),
    .B(_1079_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5493_ (.I(\as2650.pc[1] ),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5494_ (.I(_1080_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5495_ (.I(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5496_ (.A1(_3884_),
    .A2(_1008_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5497_ (.A1(_3986_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5498_ (.I(_1084_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5499_ (.I(_4081_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5500_ (.A1(_1086_),
    .A2(_1085_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5501_ (.A1(_1082_),
    .A2(_1085_),
    .B(_1087_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5502_ (.I(_1088_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5503_ (.I(_1077_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5504_ (.A1(\as2650.stack[0][1] ),
    .A2(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5505_ (.A1(_1067_),
    .A2(_1089_),
    .B(_1091_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5506_ (.I(\as2650.pc[2] ),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5507_ (.I(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5508_ (.I(_0949_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5509_ (.A1(_1094_),
    .A2(_1084_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5510_ (.A1(_1093_),
    .A2(_1085_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5511_ (.I(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5512_ (.A1(\as2650.stack[0][2] ),
    .A2(_1090_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5513_ (.A1(_1067_),
    .A2(_1097_),
    .B(_1098_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5514_ (.I(\as2650.pc[3] ),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5515_ (.I(_1099_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5516_ (.I(_0962_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5517_ (.I0(_1100_),
    .I1(_1101_),
    .S(_1074_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5518_ (.I(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5519_ (.A1(\as2650.stack[0][3] ),
    .A2(_1090_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5520_ (.A1(_1067_),
    .A2(_1103_),
    .B(_1104_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5521_ (.I(_1066_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5522_ (.I(\as2650.pc[4] ),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5523_ (.I(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5524_ (.I(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5525_ (.I(_0520_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5526_ (.I(_1013_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5527_ (.I0(_1108_),
    .I1(_1109_),
    .S(_1110_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5528_ (.I(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5529_ (.A1(\as2650.stack[0][4] ),
    .A2(_1090_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5530_ (.A1(_1105_),
    .A2(_1112_),
    .B(_1113_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5531_ (.I(\as2650.pc[5] ),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5532_ (.I(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5533_ (.I(_1115_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5534_ (.I(_0986_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5535_ (.A1(_1117_),
    .A2(_1084_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5536_ (.A1(_1116_),
    .A2(_1085_),
    .B(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5537_ (.I(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5538_ (.I(_1077_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5539_ (.A1(\as2650.stack[0][5] ),
    .A2(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5540_ (.A1(_1105_),
    .A2(_1120_),
    .B(_1122_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5541_ (.I(\as2650.pc[6] ),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5542_ (.I(_0710_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5543_ (.I(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5544_ (.I0(_1123_),
    .I1(_1125_),
    .S(_1110_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5545_ (.I(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5546_ (.A1(\as2650.stack[0][6] ),
    .A2(_1121_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5547_ (.A1(_1105_),
    .A2(_1127_),
    .B(_1128_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5548_ (.I(\as2650.pc[7] ),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5549_ (.I0(_1129_),
    .I1(_1004_),
    .S(_1110_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5550_ (.I(_1130_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5551_ (.A1(\as2650.stack[0][7] ),
    .A2(_1121_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5552_ (.A1(_1105_),
    .A2(_1131_),
    .B(_1132_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5553_ (.A1(_0884_),
    .A2(_1010_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5554_ (.A1(_1133_),
    .A2(_1064_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5555_ (.I(_1134_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5556_ (.I(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5557_ (.I(_1134_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5558_ (.I(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5559_ (.A1(\as2650.stack[1][0] ),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5560_ (.A1(_1076_),
    .A2(_1136_),
    .B(_1139_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5561_ (.I(_1137_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5562_ (.A1(\as2650.stack[1][1] ),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5563_ (.A1(_1089_),
    .A2(_1136_),
    .B(_1141_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5564_ (.A1(\as2650.stack[1][2] ),
    .A2(_1140_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5565_ (.A1(_1097_),
    .A2(_1136_),
    .B(_1142_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5566_ (.A1(\as2650.stack[1][3] ),
    .A2(_1140_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5567_ (.A1(_1103_),
    .A2(_1136_),
    .B(_1143_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5568_ (.I(_1135_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5569_ (.A1(\as2650.stack[1][4] ),
    .A2(_1140_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5570_ (.A1(_1112_),
    .A2(_1144_),
    .B(_1145_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5571_ (.I(_1137_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5572_ (.A1(\as2650.stack[1][5] ),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5573_ (.A1(_1120_),
    .A2(_1144_),
    .B(_1147_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5574_ (.A1(\as2650.stack[1][6] ),
    .A2(_1146_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5575_ (.A1(_1127_),
    .A2(_1144_),
    .B(_1148_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5576_ (.A1(\as2650.stack[1][7] ),
    .A2(_1146_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5577_ (.A1(_1131_),
    .A2(_1144_),
    .B(_1149_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5578_ (.A1(_0894_),
    .A2(_1012_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5579_ (.A1(_0887_),
    .A2(_1010_),
    .B(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5580_ (.A1(_1151_),
    .A2(_1063_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5581_ (.A1(_1011_),
    .A2(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5582_ (.I(_1153_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5583_ (.I(_1154_),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5584_ (.I(_1013_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5585_ (.I(\as2650.pc[8] ),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5586_ (.I(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5587_ (.I(_1158_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5588_ (.A1(_1159_),
    .A2(_1156_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5589_ (.A1(_4158_),
    .A2(_1156_),
    .B(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5590_ (.I(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5591_ (.I(_1154_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5592_ (.A1(\as2650.stack[2][8] ),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5593_ (.A1(_1155_),
    .A2(_1162_),
    .B(_1164_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5594_ (.I(\as2650.pc[9] ),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5595_ (.I(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5596_ (.A1(_1166_),
    .A2(_1074_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5597_ (.A1(_4260_),
    .A2(_1156_),
    .B(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5598_ (.I(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5599_ (.I(_1154_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5600_ (.A1(\as2650.stack[2][9] ),
    .A2(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5601_ (.A1(_1155_),
    .A2(_1169_),
    .B(_1171_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5602_ (.I(\as2650.pc[10] ),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5603_ (.A1(_1172_),
    .A2(_1074_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5604_ (.A1(_0369_),
    .A2(_1156_),
    .B(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5605_ (.I(_1174_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5606_ (.A1(\as2650.stack[2][10] ),
    .A2(_1170_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5607_ (.A1(_1155_),
    .A2(_1175_),
    .B(_1176_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5608_ (.I(\as2650.pc[11] ),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5609_ (.I(_1177_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5610_ (.I(_1084_),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5611_ (.A1(_0472_),
    .A2(_1110_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5612_ (.A1(_1178_),
    .A2(_1179_),
    .B(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5613_ (.I(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5614_ (.A1(\as2650.stack[2][11] ),
    .A2(_1170_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5615_ (.A1(_1155_),
    .A2(_1182_),
    .B(_1183_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5616_ (.I(\as2650.pc[12] ),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5617_ (.I(_1184_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5618_ (.I(_0568_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5619_ (.A1(_1186_),
    .A2(_1073_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5620_ (.A1(_1185_),
    .A2(_1179_),
    .B(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5621_ (.I(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5622_ (.A1(\as2650.stack[2][12] ),
    .A2(_1170_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5623_ (.A1(_1163_),
    .A2(_1189_),
    .B(_1190_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5624_ (.I(\as2650.pc[13] ),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5625_ (.A1(_0528_),
    .A2(_1073_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5626_ (.A1(_1191_),
    .A2(_1179_),
    .B(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5627_ (.I(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5628_ (.I(_1154_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5629_ (.A1(\as2650.stack[2][13] ),
    .A2(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5630_ (.A1(_1163_),
    .A2(_1194_),
    .B(_1196_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5631_ (.I(_0741_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5632_ (.A1(_1197_),
    .A2(_1073_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5633_ (.A1(\as2650.pc[14] ),
    .A2(_1179_),
    .B(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5634_ (.I(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5635_ (.A1(\as2650.stack[2][14] ),
    .A2(_1195_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5636_ (.A1(_1163_),
    .A2(_1200_),
    .B(_1201_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5637_ (.I(_1077_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5638_ (.A1(\as2650.stack[0][8] ),
    .A2(_1121_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5639_ (.A1(_1202_),
    .A2(_1162_),
    .B(_1203_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5640_ (.I(_1065_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5641_ (.A1(\as2650.stack[0][9] ),
    .A2(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5642_ (.A1(_1202_),
    .A2(_1169_),
    .B(_1205_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5643_ (.A1(\as2650.stack[0][10] ),
    .A2(_1204_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5644_ (.A1(_1202_),
    .A2(_1175_),
    .B(_1206_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5645_ (.A1(\as2650.stack[0][11] ),
    .A2(_1204_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5646_ (.A1(_1202_),
    .A2(_1182_),
    .B(_1207_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5647_ (.A1(\as2650.stack[0][12] ),
    .A2(_1204_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5648_ (.A1(_1078_),
    .A2(_1189_),
    .B(_1208_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5649_ (.A1(\as2650.stack[0][13] ),
    .A2(_1066_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5650_ (.A1(_1078_),
    .A2(_1194_),
    .B(_1209_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5651_ (.A1(\as2650.stack[0][14] ),
    .A2(_1066_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5652_ (.A1(_1078_),
    .A2(_1200_),
    .B(_1210_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5653_ (.I(_1137_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5654_ (.A1(\as2650.stack[1][8] ),
    .A2(_1146_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5655_ (.A1(_1211_),
    .A2(_1162_),
    .B(_1212_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5656_ (.I(_1134_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(\as2650.stack[1][9] ),
    .A2(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_1211_),
    .A2(_1169_),
    .B(_1214_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5659_ (.A1(\as2650.stack[1][10] ),
    .A2(_1213_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5660_ (.A1(_1211_),
    .A2(_1175_),
    .B(_1215_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5661_ (.A1(\as2650.stack[1][11] ),
    .A2(_1213_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5662_ (.A1(_1211_),
    .A2(_1182_),
    .B(_1216_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(\as2650.stack[1][12] ),
    .A2(_1213_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5664_ (.A1(_1138_),
    .A2(_1189_),
    .B(_1217_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5665_ (.A1(\as2650.stack[1][13] ),
    .A2(_1135_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5666_ (.A1(_1138_),
    .A2(_1194_),
    .B(_1218_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5667_ (.A1(\as2650.stack[1][14] ),
    .A2(_1135_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5668_ (.A1(_1138_),
    .A2(_1200_),
    .B(_1219_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5669_ (.I(\as2650.r123_2[3][0] ),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5670_ (.I(_1220_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5671_ (.I(\as2650.r123_2[3][1] ),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5672_ (.I(_1221_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5673_ (.I(\as2650.r123_2[3][2] ),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5674_ (.I(_1222_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5675_ (.I(\as2650.r123_2[3][3] ),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5676_ (.I(_1223_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5677_ (.I(\as2650.r123_2[3][4] ),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5678_ (.I(_1224_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5679_ (.I(\as2650.r123_2[3][5] ),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5680_ (.I(_1225_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5681_ (.I(\as2650.r123_2[3][6] ),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5682_ (.I(_1226_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5683_ (.I(\as2650.r123_2[3][7] ),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5684_ (.I(_1227_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5685_ (.I(_1075_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5686_ (.I(_1153_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5688_ (.A1(\as2650.stack[2][0] ),
    .A2(_1195_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5689_ (.A1(_1228_),
    .A2(_1230_),
    .B(_1231_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5690_ (.I(_1088_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5691_ (.A1(\as2650.stack[2][1] ),
    .A2(_1195_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5692_ (.A1(_1232_),
    .A2(_1230_),
    .B(_1233_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5693_ (.I(_1096_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(_1153_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5695_ (.A1(\as2650.stack[2][2] ),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5696_ (.A1(_1234_),
    .A2(_1230_),
    .B(_1236_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5697_ (.I(_1102_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5698_ (.A1(\as2650.stack[2][3] ),
    .A2(_1235_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5699_ (.A1(_1237_),
    .A2(_1230_),
    .B(_1238_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5700_ (.I(_1111_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5701_ (.I(_1229_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5702_ (.A1(\as2650.stack[2][4] ),
    .A2(_1235_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5703_ (.A1(_1239_),
    .A2(_1240_),
    .B(_1241_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5704_ (.I(_1119_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5705_ (.A1(\as2650.stack[2][5] ),
    .A2(_1235_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5706_ (.A1(_1242_),
    .A2(_1240_),
    .B(_1243_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5707_ (.I(_1126_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5708_ (.A1(\as2650.stack[2][6] ),
    .A2(_1229_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5709_ (.A1(_1244_),
    .A2(_1240_),
    .B(_1245_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5710_ (.I(_1130_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5711_ (.A1(\as2650.stack[2][7] ),
    .A2(_1229_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5712_ (.A1(_1246_),
    .A2(_1240_),
    .B(_1247_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5713_ (.A1(_1133_),
    .A2(_1152_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5714_ (.I(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5715_ (.I(_1249_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5716_ (.I(_1248_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5717_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5718_ (.A1(\as2650.stack[3][0] ),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5719_ (.A1(_1228_),
    .A2(_1250_),
    .B(_1253_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5720_ (.I(_1251_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5721_ (.A1(\as2650.stack[3][1] ),
    .A2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5722_ (.A1(_1232_),
    .A2(_1250_),
    .B(_1255_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5723_ (.A1(\as2650.stack[3][2] ),
    .A2(_1254_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5724_ (.A1(_1234_),
    .A2(_1250_),
    .B(_1256_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5725_ (.A1(\as2650.stack[3][3] ),
    .A2(_1254_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5726_ (.A1(_1237_),
    .A2(_1250_),
    .B(_1257_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5727_ (.I(_1249_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5728_ (.A1(\as2650.stack[3][4] ),
    .A2(_1254_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5729_ (.A1(_1239_),
    .A2(_1258_),
    .B(_1259_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5730_ (.I(_1251_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5731_ (.A1(\as2650.stack[3][5] ),
    .A2(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5732_ (.A1(_1242_),
    .A2(_1258_),
    .B(_1261_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5733_ (.A1(\as2650.stack[3][6] ),
    .A2(_1260_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5734_ (.A1(_1244_),
    .A2(_1258_),
    .B(_1262_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5735_ (.A1(\as2650.stack[3][7] ),
    .A2(_1260_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5736_ (.A1(_1246_),
    .A2(_1258_),
    .B(_1263_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5737_ (.A1(_1023_),
    .A2(_1061_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5738_ (.A1(_1011_),
    .A2(_1151_),
    .A3(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5739_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5740_ (.I(_1266_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5741_ (.I(_1265_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5742_ (.I(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5743_ (.A1(\as2650.stack[4][0] ),
    .A2(_1269_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5744_ (.A1(_1228_),
    .A2(_1267_),
    .B(_1270_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5745_ (.I(_1268_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5746_ (.A1(\as2650.stack[4][1] ),
    .A2(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5747_ (.A1(_1232_),
    .A2(_1267_),
    .B(_1272_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5748_ (.A1(\as2650.stack[4][2] ),
    .A2(_1271_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5749_ (.A1(_1234_),
    .A2(_1267_),
    .B(_1273_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5750_ (.A1(\as2650.stack[4][3] ),
    .A2(_1271_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5751_ (.A1(_1237_),
    .A2(_1267_),
    .B(_1274_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5752_ (.I(_1266_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5753_ (.A1(\as2650.stack[4][4] ),
    .A2(_1271_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5754_ (.A1(_1239_),
    .A2(_1275_),
    .B(_1276_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5755_ (.I(_1268_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5756_ (.A1(\as2650.stack[4][5] ),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5757_ (.A1(_1242_),
    .A2(_1275_),
    .B(_1278_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5758_ (.A1(\as2650.stack[4][6] ),
    .A2(_1277_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5759_ (.A1(_1244_),
    .A2(_1275_),
    .B(_1279_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5760_ (.A1(\as2650.stack[4][7] ),
    .A2(_1277_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5761_ (.A1(_1246_),
    .A2(_1275_),
    .B(_1280_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5762_ (.I(\as2650.psu[5] ),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5763_ (.A1(_4135_),
    .A2(_0854_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5764_ (.A1(_0461_),
    .A2(_4133_),
    .A3(_0523_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5765_ (.A1(_0847_),
    .A2(_3973_),
    .A3(_0863_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5766_ (.A1(_1008_),
    .A2(_1283_),
    .A3(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5767_ (.A1(_1282_),
    .A2(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5768_ (.A1(_3942_),
    .A2(_3914_),
    .A3(_3866_),
    .A4(_0354_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5769_ (.A1(_1287_),
    .A2(_4206_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5770_ (.A1(_3912_),
    .A2(_0850_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5771_ (.A1(_3945_),
    .A2(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5772_ (.A1(_1288_),
    .A2(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5773_ (.A1(_3884_),
    .A2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5774_ (.A1(_1286_),
    .A2(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5775_ (.I(_1289_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5776_ (.I(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5777_ (.I(_4129_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5778_ (.I(_0529_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5779_ (.A1(\as2650.psl[6] ),
    .A2(_1297_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5780_ (.I(\as2650.psl[7] ),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5781_ (.A1(_1299_),
    .A2(_0847_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5782_ (.A1(\as2650.psl[7] ),
    .A2(_0522_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5783_ (.A1(_1298_),
    .A2(_1300_),
    .A3(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5784_ (.A1(_1053_),
    .A2(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5785_ (.A1(_1296_),
    .A2(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5786_ (.I(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5787_ (.A1(_0840_),
    .A2(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5788_ (.A1(_4135_),
    .A2(_0855_),
    .A3(_1058_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5789_ (.I(_1007_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5790_ (.A1(_1308_),
    .A2(_1284_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5791_ (.A1(_1307_),
    .A2(_1309_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5792_ (.I(_1043_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5793_ (.I(_1311_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5794_ (.I(_1026_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5795_ (.I(_3879_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5796_ (.A1(_1313_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5797_ (.I(_1315_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5798_ (.I(_1316_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5799_ (.I(_1288_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5800_ (.A1(_3920_),
    .A2(_3995_),
    .A3(_3932_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5801_ (.A1(_1318_),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5802_ (.A1(_1312_),
    .A2(_1317_),
    .A3(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5803_ (.I(_1029_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5804_ (.I(_1322_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5805_ (.I(_1053_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5806_ (.I(_3983_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5807_ (.A1(_3920_),
    .A2(_3940_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5808_ (.I(_1326_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5809_ (.A1(_1325_),
    .A2(_4143_),
    .A3(_1327_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5810_ (.A1(_1324_),
    .A2(_1328_),
    .B(_1291_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5811_ (.A1(_1323_),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5812_ (.A1(_1310_),
    .A2(_1321_),
    .A3(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5813_ (.I(_3947_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5814_ (.I(_1332_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5815_ (.A1(_0530_),
    .A2(_1328_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5816_ (.I(_1027_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(_1031_),
    .A2(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5818_ (.A1(_1025_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5819_ (.A1(_3953_),
    .A2(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5820_ (.A1(_1333_),
    .A2(_1334_),
    .B(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5821_ (.A1(_1295_),
    .A2(_1306_),
    .B(_1331_),
    .C(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5822_ (.A1(_1293_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5823_ (.A1(_1052_),
    .A2(_3933_),
    .A3(_4164_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5824_ (.I(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5825_ (.I(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5826_ (.A1(_0613_),
    .A2(_0460_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5827_ (.I(_0618_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5828_ (.I(_1059_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5829_ (.I(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5830_ (.I(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5831_ (.A1(_1325_),
    .A2(_4143_),
    .A3(_1326_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5832_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5833_ (.A1(_4082_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5834_ (.A1(_1346_),
    .A2(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5835_ (.A1(\as2650.psu[5] ),
    .A2(_1346_),
    .B(_1349_),
    .C(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5836_ (.A1(_1345_),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5837_ (.A1(_1344_),
    .A2(_1355_),
    .B(_1341_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5838_ (.I(_4128_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5839_ (.I(_1357_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5840_ (.I(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5841_ (.A1(_1281_),
    .A2(_1341_),
    .B(_1356_),
    .C(_1359_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5842_ (.I(_1358_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5843_ (.I(\as2650.psl[6] ),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5844_ (.I(_3933_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5845_ (.I(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5846_ (.A1(_1031_),
    .A2(_1025_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5847_ (.I(_3875_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5848_ (.A1(_1365_),
    .A2(_1342_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5849_ (.A1(_1364_),
    .A2(_1320_),
    .A3(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5850_ (.I(_4102_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5851_ (.A1(_0444_),
    .A2(_4133_),
    .A3(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5852_ (.A1(_1286_),
    .A2(_1369_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5853_ (.A1(_3874_),
    .A2(_3932_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5854_ (.A1(_0443_),
    .A2(_4133_),
    .A3(_0530_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5855_ (.A1(_1372_),
    .A2(_1292_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5856_ (.A1(_0464_),
    .A2(_4164_),
    .A3(_1371_),
    .A4(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5857_ (.A1(_1363_),
    .A2(_1367_),
    .B1(_1370_),
    .B2(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5858_ (.I(_1048_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5859_ (.I(_1308_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5860_ (.A1(_1376_),
    .A2(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5861_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5862_ (.A1(_3967_),
    .A2(_3985_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5863_ (.A1(_0461_),
    .A2(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5864_ (.I(_1381_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5865_ (.I(_1364_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5866_ (.I(_4012_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5867_ (.A1(_1384_),
    .A2(_1319_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5868_ (.I(_3867_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5869_ (.A1(_4076_),
    .A2(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5870_ (.A1(_1385_),
    .A2(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5871_ (.I(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5872_ (.A1(_3941_),
    .A2(_1319_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5873_ (.A1(_3903_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5874_ (.I(_1308_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5875_ (.A1(_1043_),
    .A2(_3910_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5876_ (.I(_1393_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5877_ (.A1(_1392_),
    .A2(_4072_),
    .B1(_1394_),
    .B2(_4207_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5878_ (.A1(_1383_),
    .A2(_1389_),
    .B(_1391_),
    .C(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5879_ (.A1(_1379_),
    .A2(_1382_),
    .B(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5880_ (.A1(_1044_),
    .A2(_1294_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5881_ (.I(_3947_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5882_ (.A1(_1048_),
    .A2(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5883_ (.A1(_3847_),
    .A2(_1399_),
    .A3(_1350_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5884_ (.A1(_1400_),
    .A2(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5885_ (.A1(_3954_),
    .A2(_1398_),
    .A3(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5886_ (.A1(_3867_),
    .A2(_3861_),
    .A3(_3972_),
    .A4(_3918_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5887_ (.A1(_1007_),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5888_ (.A1(_1007_),
    .A2(_1283_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5889_ (.A1(_1307_),
    .A2(_1405_),
    .A3(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5890_ (.I(_1371_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5891_ (.A1(_3875_),
    .A2(_3910_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5892_ (.I(_1409_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5893_ (.I(_3946_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5894_ (.A1(_1410_),
    .A2(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5895_ (.I(_1386_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5896_ (.A1(_1413_),
    .A2(_1059_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5897_ (.A1(_1399_),
    .A2(_3963_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5898_ (.I(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5899_ (.A1(_1414_),
    .A2(_1416_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5900_ (.A1(_1412_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5901_ (.A1(_0603_),
    .A2(_1330_),
    .A3(_1408_),
    .B(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5902_ (.A1(_4021_),
    .A2(_1386_),
    .A3(_4164_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5903_ (.A1(_1420_),
    .A2(_1404_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5904_ (.A1(_1413_),
    .A2(_4129_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5905_ (.I(_1422_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5906_ (.A1(_4204_),
    .A2(_1421_),
    .A3(_1423_),
    .A4(_1382_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5907_ (.A1(_1403_),
    .A2(_1407_),
    .A3(_1419_),
    .A4(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5908_ (.A1(_1375_),
    .A2(_1397_),
    .A3(_1425_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5909_ (.A1(_1361_),
    .A2(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5910_ (.A1(_0831_),
    .A2(_0843_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5911_ (.A1(_4037_),
    .A2(_4195_),
    .A3(_0363_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5912_ (.A1(_0456_),
    .A2(_1429_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5913_ (.A1(_0510_),
    .A2(_0610_),
    .A3(_0698_),
    .A4(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5914_ (.A1(_0678_),
    .A2(_0829_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5915_ (.A1(_0587_),
    .A2(_0590_),
    .B(_1432_),
    .C(_0503_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5916_ (.I(_4130_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5917_ (.A1(_1434_),
    .A2(_4175_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5918_ (.A1(_0428_),
    .A2(_0430_),
    .B(_1435_),
    .C(_0343_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5919_ (.A1(_4008_),
    .A2(_4027_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5920_ (.A1(_1437_),
    .A2(_4175_),
    .B(_0344_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5921_ (.A1(_0343_),
    .A2(_1438_),
    .B(_0437_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5922_ (.A1(_0432_),
    .A2(_1439_),
    .B(_0504_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5923_ (.A1(_0489_),
    .A2(_0491_),
    .B1(_0503_),
    .B2(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5924_ (.A1(_0592_),
    .A2(_1441_),
    .B(_0679_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5925_ (.I(\as2650.psl[1] ),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5926_ (.A1(_0695_),
    .A2(_0685_),
    .A3(_0829_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5927_ (.A1(_1443_),
    .A2(_0830_),
    .B(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5928_ (.A1(_0826_),
    .A2(_0837_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5929_ (.I(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5930_ (.A1(_1432_),
    .A2(_1442_),
    .B(_1445_),
    .C(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5931_ (.A1(_1443_),
    .A2(_0830_),
    .A3(_1446_),
    .B(_4229_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5932_ (.I(_1392_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5933_ (.I(_1450_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5934_ (.A1(_1448_),
    .A2(_1449_),
    .B(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5935_ (.A1(_4176_),
    .A2(_1433_),
    .A3(_1436_),
    .B(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5936_ (.A1(_4229_),
    .A2(_1428_),
    .A3(_1431_),
    .B(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5937_ (.A1(_0603_),
    .A2(_1376_),
    .A3(_1325_),
    .A4(_1384_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5938_ (.I(_0825_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5939_ (.I(_1456_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5940_ (.A1(_0805_),
    .A2(_0799_),
    .B(_1455_),
    .C(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5941_ (.A1(_0290_),
    .A2(_4197_),
    .A3(_4053_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5942_ (.A1(_0710_),
    .A2(_0613_),
    .A3(_0410_),
    .A4(_0391_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5943_ (.A1(_1459_),
    .A2(_1460_),
    .B(_0817_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5944_ (.A1(_1420_),
    .A2(_1461_),
    .B(_1349_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5945_ (.I(_1376_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5946_ (.I(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5947_ (.I(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5948_ (.A1(_1458_),
    .A2(_1462_),
    .B(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5949_ (.I(_1287_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5950_ (.A1(_1467_),
    .A2(_0813_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5951_ (.A1(_1411_),
    .A2(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5952_ (.I(_1385_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5953_ (.I(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5954_ (.I(_4092_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5955_ (.I(_0413_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5956_ (.I(_0593_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5957_ (.A1(_1471_),
    .A2(_1472_),
    .A3(_1473_),
    .A4(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5958_ (.A1(_1456_),
    .A2(_0544_),
    .A3(_0690_),
    .A4(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5959_ (.I(_4207_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_1477_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5961_ (.I(_1284_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5962_ (.A1(_1479_),
    .A2(_1461_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5963_ (.A1(_1124_),
    .A2(_1479_),
    .B(_1480_),
    .C(_1450_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5964_ (.I(_1296_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5965_ (.I(_0711_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5966_ (.I(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5967_ (.I(_1484_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5968_ (.A1(_0847_),
    .A2(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5969_ (.I(_0711_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5970_ (.I(_1487_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5971_ (.I(_1488_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5972_ (.A1(_1361_),
    .A2(_1489_),
    .B(_3848_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5973_ (.A1(_1482_),
    .A2(_1351_),
    .A3(_1486_),
    .A4(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5974_ (.A1(_1478_),
    .A2(_1481_),
    .A3(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5975_ (.I(_3924_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5976_ (.I(_1493_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5977_ (.I(_1494_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5978_ (.A1(_4097_),
    .A2(_1456_),
    .B(_4024_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5979_ (.A1(_1477_),
    .A2(_0804_),
    .B(_1467_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5980_ (.A1(_1495_),
    .A2(_1496_),
    .A3(_0799_),
    .B(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5981_ (.A1(_1492_),
    .A2(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5982_ (.A1(_1469_),
    .A2(_1476_),
    .B(_1499_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5983_ (.I(_1411_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5984_ (.I(_1376_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5985_ (.I(_1502_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5986_ (.I(_1503_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5987_ (.A1(_0808_),
    .A2(_1501_),
    .B(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5988_ (.I(_1485_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5989_ (.I(_1470_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5990_ (.I(_0543_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5991_ (.I(_1508_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5992_ (.A1(_1509_),
    .A2(_0618_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5993_ (.I(_4064_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5994_ (.I(net6),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5995_ (.I(_1512_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5996_ (.I(_1513_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5997_ (.I(_1514_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5998_ (.I(_1515_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5999_ (.I(_0304_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6001_ (.I(_1518_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6002_ (.I(_0396_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6003_ (.A1(_1511_),
    .A2(_1516_),
    .A3(_1519_),
    .A4(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6004_ (.A1(_1506_),
    .A2(_1507_),
    .A3(_1510_),
    .A4(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6005_ (.A1(_1500_),
    .A2(_1505_),
    .A3(_1522_),
    .B(_1426_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6006_ (.A1(_1454_),
    .A2(_1466_),
    .B(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6007_ (.A1(_1360_),
    .A2(_1427_),
    .A3(_1524_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6008_ (.A1(_3966_),
    .A2(_0844_),
    .B(_1452_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6009_ (.A1(_0817_),
    .A2(_1434_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6010_ (.I(_1434_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6011_ (.A1(_1527_),
    .A2(_1455_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6012_ (.A1(_1457_),
    .A2(_1455_),
    .B1(_1526_),
    .B2(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6013_ (.I(_1493_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6014_ (.I(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6015_ (.I(_1482_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6016_ (.A1(_1048_),
    .A2(_4014_),
    .A3(_1326_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6017_ (.I(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6018_ (.I(_0616_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6019_ (.A1(_4016_),
    .A2(_0395_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6020_ (.A1(\as2650.psl[5] ),
    .A2(_1535_),
    .B(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6021_ (.I(\as2650.psl[7] ),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6022_ (.I(_4064_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _6023_ (.A1(_1538_),
    .A2(_0807_),
    .B1(_1539_),
    .B2(_4023_),
    .C1(\as2650.overflow ),
    .C2(_0307_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6024_ (.I(_0542_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _6025_ (.A1(\as2650.psl[1] ),
    .A2(_4225_),
    .B1(_1541_),
    .B2(_3951_),
    .C1(_1484_),
    .C2(_1361_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6026_ (.A1(_1537_),
    .A2(_1540_),
    .A3(_1542_),
    .B(_3847_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6027_ (.A1(_1534_),
    .A2(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6028_ (.I(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6029_ (.I(net3),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6030_ (.I(_1546_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6031_ (.A1(_1539_),
    .A2(_4069_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6032_ (.A1(_1547_),
    .A2(_0825_),
    .B1(_0539_),
    .B2(_0617_),
    .C(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6033_ (.I(_0713_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6034_ (.A1(_1515_),
    .A2(_4185_),
    .B1(_0312_),
    .B2(_1517_),
    .C1(_0690_),
    .C2(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6035_ (.A1(_0396_),
    .A2(_0398_),
    .B1(_0499_),
    .B2(_1508_),
    .C1(_1534_),
    .C2(_3847_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6036_ (.A1(_1549_),
    .A2(_1551_),
    .A3(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6037_ (.I(\as2650.psu[3] ),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6038_ (.A1(_0904_),
    .A2(_1517_),
    .B1(_0396_),
    .B2(_1554_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6039_ (.I(_1514_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6040_ (.A1(\as2650.psu[7] ),
    .A2(_0807_),
    .B1(_1535_),
    .B2(\as2650.psu[5] ),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _6041_ (.A1(\as2650.psu[4] ),
    .A2(_1541_),
    .B1(_1484_),
    .B2(net27),
    .C1(_0883_),
    .C2(_1539_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6042_ (.A1(_0896_),
    .A2(_1556_),
    .B(_1557_),
    .C(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6043_ (.A1(_1555_),
    .A2(_1559_),
    .B(_3848_),
    .C(_1533_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6044_ (.A1(_1368_),
    .A2(_1328_),
    .B1(_1545_),
    .B2(_1553_),
    .C(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6045_ (.I(_1546_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6046_ (.I(_1562_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6047_ (.A1(_1538_),
    .A2(_1563_),
    .A3(_1324_),
    .A4(_1351_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6048_ (.A1(_1561_),
    .A2(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6049_ (.A1(_1563_),
    .A2(_1334_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6050_ (.A1(_1334_),
    .A2(_1565_),
    .B1(_1566_),
    .B2(_1538_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6051_ (.A1(_1532_),
    .A2(_1567_),
    .B(_1526_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6052_ (.A1(_1531_),
    .A2(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6053_ (.A1(_1497_),
    .A2(_1569_),
    .B(_1469_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6054_ (.A1(_1465_),
    .A2(_1525_),
    .A3(_1529_),
    .B1(_1505_),
    .B2(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6055_ (.A1(_1538_),
    .A2(_1426_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6056_ (.A1(_1426_),
    .A2(_1571_),
    .B(_1572_),
    .C(_1359_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6057_ (.I(_1264_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6058_ (.A1(_1011_),
    .A2(_1017_),
    .A3(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6059_ (.I(_1574_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6060_ (.I(_1575_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6061_ (.I(_1574_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6062_ (.I(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6063_ (.A1(\as2650.stack[5][0] ),
    .A2(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6064_ (.A1(_1076_),
    .A2(_1576_),
    .B(_1579_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6065_ (.I(_1577_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6066_ (.A1(\as2650.stack[5][1] ),
    .A2(_1580_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6067_ (.A1(_1089_),
    .A2(_1576_),
    .B(_1581_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6068_ (.A1(\as2650.stack[5][2] ),
    .A2(_1580_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6069_ (.A1(_1097_),
    .A2(_1576_),
    .B(_1582_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6070_ (.A1(\as2650.stack[5][3] ),
    .A2(_1580_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6071_ (.A1(_1103_),
    .A2(_1576_),
    .B(_1583_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6072_ (.I(_1575_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6073_ (.A1(\as2650.stack[5][4] ),
    .A2(_1580_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6074_ (.A1(_1112_),
    .A2(_1584_),
    .B(_1585_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6075_ (.I(_1577_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6076_ (.A1(\as2650.stack[5][5] ),
    .A2(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6077_ (.A1(_1120_),
    .A2(_1584_),
    .B(_1587_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6078_ (.A1(\as2650.stack[5][6] ),
    .A2(_1586_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6079_ (.A1(_1127_),
    .A2(_1584_),
    .B(_1588_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6080_ (.A1(\as2650.stack[5][7] ),
    .A2(_1586_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6081_ (.A1(_1131_),
    .A2(_1584_),
    .B(_1589_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6082_ (.A1(_1133_),
    .A2(_1151_),
    .A3(_1573_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6083_ (.I(_1590_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6084_ (.I(_1591_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6085_ (.I(_1590_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6086_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6087_ (.A1(\as2650.stack[6][8] ),
    .A2(_1594_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6088_ (.A1(_1162_),
    .A2(_1592_),
    .B(_1595_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6089_ (.I(_1593_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6090_ (.A1(\as2650.stack[6][9] ),
    .A2(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6091_ (.A1(_1169_),
    .A2(_1592_),
    .B(_1597_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6092_ (.A1(\as2650.stack[6][10] ),
    .A2(_1596_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6093_ (.A1(_1175_),
    .A2(_1592_),
    .B(_1598_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6094_ (.A1(\as2650.stack[6][11] ),
    .A2(_1596_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6095_ (.A1(_1182_),
    .A2(_1592_),
    .B(_1599_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6096_ (.I(_1591_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6097_ (.A1(\as2650.stack[6][12] ),
    .A2(_1596_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6098_ (.A1(_1189_),
    .A2(_1600_),
    .B(_1601_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6099_ (.I(_1593_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6100_ (.A1(\as2650.stack[6][13] ),
    .A2(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6101_ (.A1(_1194_),
    .A2(_1600_),
    .B(_1603_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6102_ (.A1(\as2650.stack[6][14] ),
    .A2(_1602_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6103_ (.A1(_1200_),
    .A2(_1600_),
    .B(_1604_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6104_ (.I(_1377_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6105_ (.I(_1605_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6106_ (.I(_1315_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6107_ (.A1(_1314_),
    .A2(_3897_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6108_ (.I(_1608_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6109_ (.A1(_1052_),
    .A2(_1045_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6110_ (.I(_1610_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6111_ (.I(_1611_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6112_ (.A1(_1607_),
    .A2(_1609_),
    .A3(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6113_ (.I(_1055_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6114_ (.A1(_1024_),
    .A2(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6115_ (.I(_1615_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6116_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6117_ (.A1(_1562_),
    .A2(_1332_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6118_ (.A1(_1609_),
    .A2(_1617_),
    .B(_1618_),
    .C(_4139_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6119_ (.A1(_1606_),
    .A2(_1613_),
    .A3(_1619_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6120_ (.I(_1620_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6121_ (.I(_1511_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6122_ (.A1(_1622_),
    .A2(_1337_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6123_ (.A1(_3849_),
    .A2(_1620_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6124_ (.I(_1054_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6125_ (.A1(_1625_),
    .A2(_1337_),
    .A3(_1620_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6126_ (.A1(_1621_),
    .A2(_1623_),
    .B(_1624_),
    .C(_1626_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6127_ (.A1(_0849_),
    .A2(_1621_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6128_ (.I(_1516_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6129_ (.A1(_4139_),
    .A2(_1609_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6130_ (.I(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6131_ (.A1(_1628_),
    .A2(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6132_ (.A1(_1626_),
    .A2(_1627_),
    .A3(_1631_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6133_ (.I(_1629_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6134_ (.I(_1052_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6135_ (.I(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6136_ (.A1(_1634_),
    .A2(_1629_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6137_ (.A1(_0308_),
    .A2(_1632_),
    .B(_1635_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6138_ (.I(_1617_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6139_ (.A1(_0840_),
    .A2(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6140_ (.A1(_0840_),
    .A2(_1620_),
    .B1(_1629_),
    .B2(_1346_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6141_ (.A1(_1626_),
    .A2(_1637_),
    .B(_1638_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6142_ (.I(_1550_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6143_ (.A1(_1325_),
    .A2(_1621_),
    .B1(_1632_),
    .B2(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6144_ (.I(_1640_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6145_ (.I(_1563_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6146_ (.A1(_1384_),
    .A2(_1621_),
    .B1(_1630_),
    .B2(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6147_ (.I(_1642_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6148_ (.I(\as2650.r123[3][0] ),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6149_ (.I(_1643_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(\as2650.r123[3][1] ),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6151_ (.I(_1644_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6152_ (.I(\as2650.r123[3][2] ),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6153_ (.I(_1645_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6154_ (.I(\as2650.r123[3][3] ),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6155_ (.I(_1646_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6156_ (.I(\as2650.r123[3][4] ),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6157_ (.I(_1647_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6158_ (.I(\as2650.r123[3][5] ),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6159_ (.I(_1648_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6160_ (.I(\as2650.r123[3][6] ),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6161_ (.I(_1649_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6162_ (.I(\as2650.r123[3][7] ),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6163_ (.I(_1650_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6164_ (.A1(_3951_),
    .A2(_3850_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6165_ (.I(_1651_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6166_ (.A1(_1347_),
    .A2(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6167_ (.A1(_0464_),
    .A2(_1653_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6168_ (.I(_1654_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6169_ (.I(_1655_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6170_ (.A1(_4137_),
    .A2(_1652_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6171_ (.I(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6172_ (.A1(_3967_),
    .A2(_1651_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6173_ (.A1(_0458_),
    .A2(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6174_ (.A1(_4057_),
    .A2(_1660_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6175_ (.I(_1661_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6176_ (.I(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6177_ (.A1(_3951_),
    .A2(_3850_),
    .A3(_4082_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6178_ (.A1(_3883_),
    .A2(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6179_ (.A1(_4072_),
    .A2(_1665_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6180_ (.I(_1666_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6181_ (.I(_1667_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6182_ (.A1(_4145_),
    .A2(_1659_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6183_ (.I(_1669_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6184_ (.I(_1670_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6185_ (.A1(_1313_),
    .A2(_1335_),
    .A3(_3904_),
    .A4(_1032_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6186_ (.I(_1659_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6187_ (.A1(_1365_),
    .A2(_1385_),
    .A3(_1672_),
    .A4(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6188_ (.A1(_4070_),
    .A2(_1674_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6189_ (.I(_1666_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6190_ (.A1(_4065_),
    .A2(_1671_),
    .B(_1675_),
    .C(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6191_ (.A1(_3875_),
    .A2(_4206_),
    .A3(_1665_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6192_ (.I(_1678_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6193_ (.I(_1679_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6194_ (.A1(_0291_),
    .A2(_1668_),
    .B(_1677_),
    .C(_1680_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6195_ (.A1(_1043_),
    .A2(_1493_),
    .A3(_1660_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6196_ (.I(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6197_ (.I(_1661_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6198_ (.A1(_4111_),
    .A2(_1683_),
    .B(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6199_ (.A1(_3938_),
    .A2(_1664_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6200_ (.I(_1686_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6201_ (.A1(_4054_),
    .A2(_1663_),
    .B1(_1681_),
    .B2(_1685_),
    .C(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6202_ (.A1(_4141_),
    .A2(_1673_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6203_ (.I(_1689_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6204_ (.I(_1673_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6205_ (.A1(_4050_),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6206_ (.A1(_4047_),
    .A2(_1690_),
    .B(_1692_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6207_ (.A1(_1688_),
    .A2(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6208_ (.I(_1657_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6209_ (.A1(_4050_),
    .A2(_1673_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6210_ (.I(_1696_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6211_ (.A1(_4124_),
    .A2(_1697_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6212_ (.A1(_1695_),
    .A2(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6213_ (.A1(_4037_),
    .A2(_1658_),
    .B1(_1694_),
    .B2(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6214_ (.A1(_1656_),
    .A2(_1700_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6215_ (.A1(_3902_),
    .A2(_1664_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6216_ (.A1(_1679_),
    .A2(_1667_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6217_ (.I(_1657_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6218_ (.A1(_3985_),
    .A2(_1665_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6219_ (.I(_1705_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6220_ (.I(_3931_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6221_ (.I(_1707_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6222_ (.A1(_4140_),
    .A2(_1708_),
    .A3(_3937_),
    .A4(_1691_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6223_ (.A1(_1704_),
    .A2(_1706_),
    .A3(_1674_),
    .A4(_1709_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6224_ (.A1(_1702_),
    .A2(_1703_),
    .A3(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6225_ (.A1(_1324_),
    .A2(_1711_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6226_ (.I(_1712_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6227_ (.A1(_1687_),
    .A2(_1684_),
    .A3(_1702_),
    .A4(_1703_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6228_ (.A1(_1704_),
    .A2(_1671_),
    .A3(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6229_ (.A1(_1368_),
    .A2(_1715_),
    .B(_1654_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6230_ (.I(_1716_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6231_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_1655_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_0767_),
    .A2(_0795_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6234_ (.A1(_0767_),
    .A2(_0795_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6235_ (.A1(_0765_),
    .A2(_1720_),
    .B(_1721_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6236_ (.A1(_0773_),
    .A2(_0793_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6237_ (.A1(_0770_),
    .A2(_0794_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6238_ (.A1(_1723_),
    .A2(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6239_ (.A1(_0627_),
    .A2(_4259_),
    .A3(_0776_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6240_ (.A1(_0778_),
    .A2(_0779_),
    .B(_1726_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6241_ (.A1(_0746_),
    .A2(_0750_),
    .A3(_0791_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6242_ (.A1(_0780_),
    .A2(_0792_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6243_ (.A1(_1728_),
    .A2(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6244_ (.A1(_0408_),
    .A2(_0566_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6245_ (.A1(_0774_),
    .A2(_0783_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6246_ (.A1(_0749_),
    .A2(_1731_),
    .B1(_1732_),
    .B2(_0782_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6247_ (.A1(\as2650.r0[7] ),
    .A2(_4256_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6248_ (.A1(_1733_),
    .A2(_1734_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6249_ (.A1(_0745_),
    .A2(_0790_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6250_ (.A1(_0745_),
    .A2(_0790_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6251_ (.A1(_0784_),
    .A2(_1736_),
    .B(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6252_ (.A1(\as2650.r0[6] ),
    .A2(_0368_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6253_ (.A1(\as2650.r0[5] ),
    .A2(_0468_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6254_ (.A1(_1731_),
    .A2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6255_ (.A1(_1739_),
    .A2(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6256_ (.A1(\as2650.r0[1] ),
    .A2(_0787_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6257_ (.A1(_3999_),
    .A2(_0788_),
    .B1(_0744_),
    .B2(_0561_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6258_ (.A1(_0742_),
    .A2(_1743_),
    .B1(_1744_),
    .B2(_0786_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6259_ (.A1(\as2650.r0[3] ),
    .A2(_0525_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6260_ (.A1(_4212_),
    .A2(_0740_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6261_ (.A1(_1743_),
    .A2(_1746_),
    .A3(_1747_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6262_ (.A1(_1745_),
    .A2(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6263_ (.A1(_1742_),
    .A2(_1749_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6264_ (.A1(_1738_),
    .A2(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6265_ (.A1(_1735_),
    .A2(_1751_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6266_ (.A1(_1730_),
    .A2(_1752_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6267_ (.A1(_1727_),
    .A2(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6268_ (.A1(_1725_),
    .A2(_1754_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6269_ (.A1(_1722_),
    .A2(_1755_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6270_ (.A1(_1719_),
    .A2(_1756_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6271_ (.A1(_1701_),
    .A2(_1713_),
    .B(_1718_),
    .C(_1757_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6272_ (.I(_1704_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6273_ (.I(_1692_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6274_ (.A1(_3901_),
    .A2(_1691_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6275_ (.I(_1678_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6276_ (.I(_1666_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6277_ (.I(_4234_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6278_ (.A1(_1763_),
    .A2(_1669_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6279_ (.A1(_1556_),
    .A2(_1670_),
    .B(_1764_),
    .C(_1667_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6280_ (.A1(_0392_),
    .A2(_1762_),
    .B(_1765_),
    .C(_1679_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6281_ (.A1(_4202_),
    .A2(_1761_),
    .B(_1766_),
    .C(_1705_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6282_ (.A1(_1086_),
    .A2(_1706_),
    .B(_1767_),
    .C(_1690_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6283_ (.A1(_4245_),
    .A2(_1690_),
    .B(_1760_),
    .C(_1768_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6284_ (.A1(_4249_),
    .A2(_1759_),
    .B(_1769_),
    .C(_1704_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6285_ (.A1(_4195_),
    .A2(_1758_),
    .B(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6286_ (.A1(_1656_),
    .A2(_1771_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6287_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_1717_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6288_ (.I(_1725_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6289_ (.A1(_1722_),
    .A2(_1755_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6290_ (.A1(_1774_),
    .A2(_1754_),
    .B(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6291_ (.A1(_1730_),
    .A2(_1752_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6292_ (.A1(_1727_),
    .A2(_1753_),
    .B(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6293_ (.A1(_0816_),
    .A2(_4260_),
    .A3(_1733_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6294_ (.A1(_1738_),
    .A2(_1750_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6295_ (.A1(_1735_),
    .A2(_1751_),
    .B(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6296_ (.A1(_0532_),
    .A2(_0568_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6297_ (.A1(_0783_),
    .A2(_1782_),
    .B1(_1741_),
    .B2(_1739_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6298_ (.I(_1748_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6299_ (.A1(_1745_),
    .A2(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6300_ (.A1(_1742_),
    .A2(_1749_),
    .B(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6301_ (.A1(\as2650.r0[7] ),
    .A2(_0368_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6302_ (.A1(_0625_),
    .A2(_0471_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6303_ (.A1(_1782_),
    .A2(_1787_),
    .A3(_1788_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6304_ (.A1(_1743_),
    .A2(_1747_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6305_ (.A1(_4212_),
    .A2(_0788_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6306_ (.A1(_0785_),
    .A2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6307_ (.A1(_1746_),
    .A2(_1790_),
    .B(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6308_ (.A1(_0292_),
    .A2(_0744_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6309_ (.A1(_1791_),
    .A2(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6310_ (.A1(_0408_),
    .A2(_0526_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6311_ (.A1(_1795_),
    .A2(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6312_ (.A1(_1793_),
    .A2(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6313_ (.A1(_1789_),
    .A2(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6314_ (.A1(_1786_),
    .A2(_1799_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6315_ (.A1(_1783_),
    .A2(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6316_ (.A1(_1781_),
    .A2(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6317_ (.A1(_1779_),
    .A2(_1802_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6318_ (.A1(_1776_),
    .A2(_1778_),
    .A3(_1803_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6319_ (.A1(_1719_),
    .A2(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6320_ (.A1(_1713_),
    .A2(_1772_),
    .B(_1773_),
    .C(_1805_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6321_ (.I(_1712_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6322_ (.A1(_0464_),
    .A2(_1653_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6323_ (.I(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6324_ (.I(_1696_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6325_ (.I(_1686_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6326_ (.A1(_3948_),
    .A2(_1659_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6327_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6328_ (.A1(_4072_),
    .A2(_1665_),
    .B1(_1811_),
    .B2(_0307_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6329_ (.A1(_0318_),
    .A2(_1812_),
    .B(_1813_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6330_ (.A1(_0398_),
    .A2(_1676_),
    .B(_1814_),
    .C(_1761_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6331_ (.A1(_0291_),
    .A2(_1682_),
    .B(_1661_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6332_ (.A1(_0290_),
    .A2(_1662_),
    .B1(_1815_),
    .B2(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6333_ (.A1(_1687_),
    .A2(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6334_ (.A1(_0331_),
    .A2(_1810_),
    .B(_1697_),
    .C(_1818_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6335_ (.A1(_0337_),
    .A2(_1809_),
    .B(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6336_ (.I0(_0363_),
    .I1(_1820_),
    .S(_1695_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6337_ (.A1(_1808_),
    .A2(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6338_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_1717_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6339_ (.A1(_1786_),
    .A2(_1799_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6340_ (.A1(_1783_),
    .A2(_1800_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6341_ (.I(_1787_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6342_ (.A1(_1782_),
    .A2(_1788_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6343_ (.A1(_1782_),
    .A2(_1788_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6344_ (.A1(_1826_),
    .A2(_1827_),
    .B(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6345_ (.A1(_1793_),
    .A2(_1797_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6346_ (.A1(_1789_),
    .A2(_1798_),
    .B(_1830_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6347_ (.A1(_4098_),
    .A2(_0472_),
    .B1(_1186_),
    .B2(_0626_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6348_ (.A1(_4098_),
    .A2(_0568_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6349_ (.A1(_1788_),
    .A2(_1833_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6350_ (.I(_1834_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6351_ (.A1(_1832_),
    .A2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6352_ (.I(_0788_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6353_ (.A1(_0293_),
    .A2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6354_ (.A1(_1747_),
    .A2(_1838_),
    .B1(_1795_),
    .B2(_1796_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6355_ (.A1(_0409_),
    .A2(_0741_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6356_ (.A1(_1838_),
    .A2(_1840_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6357_ (.A1(_0533_),
    .A2(_0527_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6358_ (.A1(_1841_),
    .A2(_1842_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6359_ (.A1(_1839_),
    .A2(_1843_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6360_ (.A1(_1836_),
    .A2(_1844_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6361_ (.A1(_1831_),
    .A2(_1845_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6362_ (.A1(_1829_),
    .A2(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6363_ (.A1(_1824_),
    .A2(_1825_),
    .B(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6364_ (.A1(_1824_),
    .A2(_1825_),
    .A3(_1847_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6365_ (.A1(_1848_),
    .A2(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6366_ (.A1(_1781_),
    .A2(_1801_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6367_ (.A1(_1779_),
    .A2(_1802_),
    .B(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6368_ (.A1(_1850_),
    .A2(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6369_ (.A1(_1778_),
    .A2(_1803_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6370_ (.A1(_1778_),
    .A2(_1803_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6371_ (.A1(_1776_),
    .A2(_1854_),
    .B(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6372_ (.A1(_1853_),
    .A2(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6373_ (.A1(_1719_),
    .A2(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6374_ (.A1(_1806_),
    .A2(_1822_),
    .B(_1823_),
    .C(_1858_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6375_ (.I(_1807_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6376_ (.I(_1686_),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6377_ (.I(_1669_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6378_ (.A1(_0401_),
    .A2(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6379_ (.A1(_1520_),
    .A2(_1671_),
    .B(_1862_),
    .C(_1676_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6380_ (.A1(_0614_),
    .A2(_1668_),
    .B(_1863_),
    .C(_1680_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6381_ (.A1(_0392_),
    .A2(_1683_),
    .B(_1684_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6382_ (.A1(_0391_),
    .A2(_1663_),
    .B1(_1864_),
    .B2(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6383_ (.A1(_0422_),
    .A2(_1687_),
    .B(_1697_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6384_ (.A1(_1860_),
    .A2(_1866_),
    .B(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6385_ (.A1(_0390_),
    .A2(_1759_),
    .B(_1868_),
    .C(_1658_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6386_ (.A1(_0456_),
    .A2(_1758_),
    .B(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6387_ (.A1(_1859_),
    .A2(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6388_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_1717_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6389_ (.A1(_1850_),
    .A2(_1852_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6390_ (.A1(_1853_),
    .A2(_1856_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6391_ (.A1(_1873_),
    .A2(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6392_ (.A1(_1839_),
    .A2(_1843_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6393_ (.A1(_1836_),
    .A2(_1844_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6394_ (.A1(_1876_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6395_ (.A1(_0410_),
    .A2(_1837_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6396_ (.A1(_1794_),
    .A2(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6397_ (.A1(_1841_),
    .A2(_1842_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6398_ (.A1(_1880_),
    .A2(_1881_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6399_ (.A1(_0533_),
    .A2(_0741_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6400_ (.A1(_1879_),
    .A2(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6401_ (.A1(_0626_),
    .A2(_0527_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6402_ (.A1(_1884_),
    .A2(_1885_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6403_ (.A1(_1882_),
    .A2(_1886_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6404_ (.A1(_1833_),
    .A2(_1887_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6405_ (.A1(_1878_),
    .A2(_1888_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6406_ (.A1(_1834_),
    .A2(_1889_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6407_ (.I(_1846_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6408_ (.A1(_1831_),
    .A2(_1845_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6409_ (.A1(_1829_),
    .A2(_1891_),
    .B(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6410_ (.A1(_1890_),
    .A2(_1893_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6411_ (.A1(_1848_),
    .A2(_1875_),
    .A3(_1894_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6412_ (.A1(_1719_),
    .A2(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6413_ (.A1(_1806_),
    .A2(_1871_),
    .B(_1872_),
    .C(_1896_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6414_ (.A1(_0547_),
    .A2(_1861_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6415_ (.A1(_1508_),
    .A2(_1861_),
    .B(_1897_),
    .C(_1762_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6416_ (.A1(_0540_),
    .A2(_1668_),
    .B(_1898_),
    .C(_1680_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6417_ (.I(_0398_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6418_ (.A1(_1900_),
    .A2(_1683_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6419_ (.A1(_1899_),
    .A2(_1901_),
    .B(_1684_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6420_ (.A1(_1109_),
    .A2(_1663_),
    .B(_1902_),
    .C(_1860_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6421_ (.A1(_0518_),
    .A2(_1810_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6422_ (.A1(_1760_),
    .A2(_1904_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6423_ (.A1(_0557_),
    .A2(_1759_),
    .B1(_1903_),
    .B2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6424_ (.A1(_0511_),
    .A2(_1658_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6425_ (.A1(_1758_),
    .A2(_1906_),
    .B(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6426_ (.A1(_1859_),
    .A2(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6427_ (.I(_1716_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6428_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6429_ (.I(_1655_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6430_ (.A1(_1848_),
    .A2(_1894_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6431_ (.A1(_1848_),
    .A2(_1873_),
    .B(_1894_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6432_ (.A1(_1853_),
    .A2(_1856_),
    .A3(_1913_),
    .B(_1914_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6433_ (.A1(_1890_),
    .A2(_1893_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6434_ (.A1(_0612_),
    .A2(_1837_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6435_ (.A1(_1840_),
    .A2(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6436_ (.A1(_1884_),
    .A2(_1885_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6437_ (.A1(_1918_),
    .A2(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6438_ (.A1(_0626_),
    .A2(_1197_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6439_ (.I(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6440_ (.A1(_1917_),
    .A2(_1922_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6441_ (.A1(_4099_),
    .A2(_0528_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6442_ (.A1(_1923_),
    .A2(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6443_ (.A1(_1920_),
    .A2(_1925_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6444_ (.A1(_1920_),
    .A2(_1925_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6445_ (.A1(_1926_),
    .A2(_1927_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6446_ (.A1(_0816_),
    .A2(_1186_),
    .A3(_1887_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6447_ (.A1(_1882_),
    .A2(_1886_),
    .B(_1929_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6448_ (.A1(_1928_),
    .A2(_1930_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6449_ (.I(_1888_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6450_ (.A1(_1878_),
    .A2(_1932_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6451_ (.A1(_1834_),
    .A2(_1889_),
    .Z(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6452_ (.A1(_1933_),
    .A2(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6453_ (.A1(_1931_),
    .A2(_1935_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6454_ (.A1(_1916_),
    .A2(_1936_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6455_ (.A1(_1915_),
    .A2(_1937_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6456_ (.A1(_1912_),
    .A2(_1938_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6457_ (.A1(_1806_),
    .A2(_1909_),
    .B(_1911_),
    .C(_1939_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6458_ (.I(_0646_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6459_ (.A1(_0617_),
    .A2(_1812_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6460_ (.A1(_0622_),
    .A2(_1812_),
    .B(_1941_),
    .C(_1762_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6461_ (.A1(_0804_),
    .A2(_1668_),
    .B(_1942_),
    .C(_1761_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6462_ (.A1(_0614_),
    .A2(_1680_),
    .B(_1943_),
    .C(_1706_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6463_ (.A1(_0986_),
    .A2(_1706_),
    .B(_1944_),
    .C(_1690_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6464_ (.A1(_3901_),
    .A2(_1691_),
    .B1(_1860_),
    .B2(_0643_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6465_ (.A1(_1940_),
    .A2(_1809_),
    .B1(_1945_),
    .B2(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6466_ (.I0(_0611_),
    .I1(_1947_),
    .S(_1658_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6467_ (.A1(_1808_),
    .A2(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6468_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_1910_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6469_ (.A1(_1916_),
    .A2(_1936_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6470_ (.A1(_1915_),
    .A2(_1937_),
    .B(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6471_ (.A1(_1933_),
    .A2(_1934_),
    .B(_1931_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6472_ (.I(_1928_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6473_ (.A1(_1954_),
    .A2(_1930_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6474_ (.A1(_1926_),
    .A2(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6475_ (.I(_1837_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6476_ (.A1(_0627_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6477_ (.A1(_1883_),
    .A2(_1958_),
    .B1(_1923_),
    .B2(_1924_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6478_ (.A1(_4099_),
    .A2(_1197_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6479_ (.A1(_1958_),
    .A2(_1960_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6480_ (.A1(_1959_),
    .A2(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6481_ (.A1(_1956_),
    .A2(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6482_ (.A1(_1953_),
    .A2(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6483_ (.A1(_1952_),
    .A2(_1964_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6484_ (.A1(_1912_),
    .A2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6485_ (.A1(_1806_),
    .A2(_1949_),
    .B(_1950_),
    .C(_1966_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6486_ (.A1(_1953_),
    .A2(_1963_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6487_ (.A1(_1952_),
    .A2(_1964_),
    .B(_1967_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6488_ (.A1(_1955_),
    .A2(_1962_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6489_ (.A1(_0816_),
    .A2(_1957_),
    .A3(_1921_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6490_ (.A1(_1959_),
    .A2(_1961_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6491_ (.A1(_1926_),
    .A2(_1962_),
    .B(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6492_ (.A1(_1970_),
    .A2(_1972_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6493_ (.A1(_1969_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6494_ (.A1(_1968_),
    .A2(_1974_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6495_ (.I(_0698_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6496_ (.A1(_0998_),
    .A2(_1662_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6497_ (.A1(_0718_),
    .A2(_1670_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6498_ (.A1(_1550_),
    .A2(_1670_),
    .B(_1978_),
    .C(_1667_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6499_ (.A1(_0825_),
    .A2(_1762_),
    .B(_1979_),
    .C(_1679_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6500_ (.A1(_1474_),
    .A2(_1761_),
    .B(_1980_),
    .C(_1705_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6501_ (.A1(_1977_),
    .A2(_1981_),
    .B(_1686_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6502_ (.A1(_0709_),
    .A2(_1810_),
    .B(_1697_),
    .C(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6503_ (.A1(_0706_),
    .A2(_1809_),
    .B(_1983_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6504_ (.I0(_1976_),
    .I1(_1984_),
    .S(_1695_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6505_ (.A1(_1808_),
    .A2(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6506_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_1910_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6507_ (.A1(_1859_),
    .A2(_1975_),
    .B1(_1986_),
    .B2(_1713_),
    .C(_1987_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6508_ (.A1(_1922_),
    .A2(_1972_),
    .B(_1957_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6509_ (.A1(_1955_),
    .A2(_1962_),
    .A3(_1973_),
    .B1(_1988_),
    .B2(_1004_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6510_ (.A1(_1968_),
    .A2(_1974_),
    .B(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6511_ (.A1(_0810_),
    .A2(_1861_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6512_ (.A1(_0807_),
    .A2(_1671_),
    .B(_1991_),
    .C(_1676_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6513_ (.A1(_0813_),
    .A2(_1682_),
    .B(_1703_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6514_ (.A1(_0804_),
    .A2(_1683_),
    .B1(_1992_),
    .B2(_1993_),
    .C(_1662_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6515_ (.A1(_1003_),
    .A2(_1663_),
    .B(_1994_),
    .C(_1810_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6516_ (.A1(_0803_),
    .A2(_1860_),
    .B(_1809_),
    .C(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6517_ (.A1(_0822_),
    .A2(_1759_),
    .B(_1695_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6518_ (.A1(_0844_),
    .A2(_1758_),
    .B1(_1996_),
    .B2(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6519_ (.A1(_1808_),
    .A2(_1998_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6520_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_1910_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6521_ (.A1(_1859_),
    .A2(_1990_),
    .B1(_1999_),
    .B2(_1713_),
    .C(_2000_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6522_ (.A1(_3849_),
    .A2(_1711_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6523_ (.I(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6524_ (.I(_1812_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6525_ (.A1(_1657_),
    .A2(_1689_),
    .A3(_1705_),
    .A4(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6526_ (.A1(_2004_),
    .A2(_1702_),
    .A3(_1703_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6527_ (.A1(_3849_),
    .A2(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6528_ (.A1(_1655_),
    .A2(_2006_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6529_ (.I(_2007_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6530_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6531_ (.A1(_4153_),
    .A2(_4158_),
    .A3(_1912_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6532_ (.A1(_1701_),
    .A2(_2002_),
    .B(_2009_),
    .C(_2010_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6533_ (.I(_2001_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6534_ (.A1(_0287_),
    .A2(_1656_),
    .B1(_2008_),
    .B2(\as2650.r123_2[1][1] ),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6535_ (.A1(_1772_),
    .A2(_2011_),
    .B(_2012_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6536_ (.A1(\as2650.r123_2[1][2] ),
    .A2(_2008_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6537_ (.A1(_0375_),
    .A2(_1912_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6538_ (.A1(_1822_),
    .A2(_2002_),
    .B(_2013_),
    .C(_2014_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6539_ (.I(_2007_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6540_ (.I(_1807_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6541_ (.A1(_0482_),
    .A2(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6542_ (.A1(\as2650.r123_2[1][3] ),
    .A2(_2015_),
    .B(_2017_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6543_ (.A1(_1871_),
    .A2(_2011_),
    .B(_2018_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6544_ (.A1(_0584_),
    .A2(_1656_),
    .B1(_2008_),
    .B2(\as2650.r123_2[1][4] ),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6545_ (.A1(_1909_),
    .A2(_2011_),
    .B(_2019_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6546_ (.A1(_0673_),
    .A2(_2016_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6547_ (.A1(\as2650.r123_2[1][5] ),
    .A2(_2015_),
    .B(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6548_ (.A1(_1949_),
    .A2(_2011_),
    .B(_2021_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6549_ (.A1(_0761_),
    .A2(_2016_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6550_ (.A1(\as2650.r123_2[1][6] ),
    .A2(_2015_),
    .B(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6551_ (.A1(_1986_),
    .A2(_2002_),
    .B(_2023_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6552_ (.A1(_0796_),
    .A2(_2016_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6553_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_2015_),
    .B(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6554_ (.A1(_1999_),
    .A2(_2002_),
    .B(_2025_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6555_ (.A1(_0848_),
    .A2(_2005_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6556_ (.I(_2026_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6557_ (.I(_2026_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6558_ (.A1(_1606_),
    .A2(_0856_),
    .A3(_1652_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6559_ (.I(_2029_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6560_ (.A1(_0458_),
    .A2(_0851_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6561_ (.A1(_2031_),
    .A2(_1652_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6562_ (.I(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6563_ (.I(_2029_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6564_ (.A1(_0865_),
    .A2(_0912_),
    .B1(_2033_),
    .B2(_1072_),
    .C(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6565_ (.A1(\as2650.r123_2[0][0] ),
    .A2(_2028_),
    .A3(_2030_),
    .B(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6566_ (.A1(_1700_),
    .A2(_2027_),
    .B(_2036_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6567_ (.I(_1372_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6568_ (.A1(_0864_),
    .A2(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6569_ (.A1(_2038_),
    .A2(_1653_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6570_ (.I(_2039_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6571_ (.A1(_1771_),
    .A2(_2026_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6572_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_2027_),
    .B(_2040_),
    .C(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6573_ (.A1(_4198_),
    .A2(_2033_),
    .B(_2030_),
    .C(_0928_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6574_ (.A1(_2042_),
    .A2(_2043_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6575_ (.A1(_0848_),
    .A2(_2005_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6576_ (.I(_2044_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6577_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_2045_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6578_ (.A1(_1821_),
    .A2(_2027_),
    .B(_2030_),
    .C(_2046_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6579_ (.A1(_0871_),
    .A2(_1653_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6580_ (.A1(_0948_),
    .A2(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6581_ (.A1(_0949_),
    .A2(_2032_),
    .B(_2049_),
    .C(_2040_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6582_ (.A1(_2047_),
    .A2(_2050_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6583_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_2045_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6584_ (.A1(_1870_),
    .A2(_2028_),
    .B(_2034_),
    .C(_2051_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6585_ (.I(_0961_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6586_ (.I(_2039_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6587_ (.A1(_0962_),
    .A2(_0865_),
    .B1(_2053_),
    .B2(_2033_),
    .C(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6588_ (.A1(_2052_),
    .A2(_2055_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6589_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_2044_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6590_ (.A1(_1908_),
    .A2(_2028_),
    .B(_2034_),
    .C(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6591_ (.A1(_0973_),
    .A2(_2048_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6592_ (.A1(_0519_),
    .A2(_2032_),
    .B(_2058_),
    .C(_2054_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6593_ (.A1(_2057_),
    .A2(_2059_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6594_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_2044_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6595_ (.A1(_1948_),
    .A2(_2028_),
    .B(_2034_),
    .C(_2060_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6596_ (.I(_0985_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6597_ (.A1(_0967_),
    .A2(_2062_),
    .B1(_2048_),
    .B2(_0986_),
    .C(_2054_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6598_ (.A1(_2061_),
    .A2(_2063_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6599_ (.A1(\as2650.r123_2[0][6] ),
    .A2(_2045_),
    .B(_2030_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6600_ (.A1(_1985_),
    .A2(_2027_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6601_ (.A1(_0997_),
    .A2(_2048_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6602_ (.A1(_0998_),
    .A2(_2032_),
    .B(_2066_),
    .C(_2054_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6603_ (.A1(_2064_),
    .A2(_2065_),
    .B(_2067_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6604_ (.I(_1004_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6605_ (.A1(\as2650.r123_2[0][7] ),
    .A2(_2026_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6606_ (.A1(_1998_),
    .A2(_2045_),
    .B(_2040_),
    .C(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6607_ (.A1(_2068_),
    .A2(_0967_),
    .A3(_2040_),
    .B(_2070_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6608_ (.I(_1539_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6609_ (.A1(_3895_),
    .A2(_3881_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6610_ (.I(_2072_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6611_ (.A1(_1314_),
    .A2(_2073_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6612_ (.I(_3890_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6613_ (.A1(\as2650.cycle[7] ),
    .A2(_3929_),
    .A3(_2072_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6614_ (.I(_2076_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6615_ (.A1(_2075_),
    .A2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6616_ (.A1(_1413_),
    .A2(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6617_ (.A1(_2074_),
    .A2(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6618_ (.A1(_3958_),
    .A2(_1039_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6619_ (.A1(_4048_),
    .A2(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6620_ (.A1(_1026_),
    .A2(_1335_),
    .A3(_3904_),
    .A4(_1032_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6621_ (.A1(_1024_),
    .A2(_1045_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6622_ (.I(_2084_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6623_ (.A1(_2083_),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6624_ (.A1(_3962_),
    .A2(_2086_),
    .B(_3955_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6625_ (.A1(_2080_),
    .A2(_2082_),
    .A3(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6626_ (.I(_1034_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6627_ (.A1(_1386_),
    .A2(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6628_ (.I(_2090_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6629_ (.A1(_1337_),
    .A2(_1400_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6630_ (.A1(_3954_),
    .A2(_2091_),
    .A3(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6631_ (.A1(_1029_),
    .A2(_1034_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6632_ (.A1(_1044_),
    .A2(_1057_),
    .A3(_2094_),
    .A4(_2081_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6633_ (.A1(_1377_),
    .A2(_1040_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6634_ (.I(_1413_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6635_ (.A1(_1707_),
    .A2(_2096_),
    .B(_2097_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6636_ (.A1(_4130_),
    .A2(_2095_),
    .B(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6637_ (.A1(_2093_),
    .A2(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6638_ (.I(_2089_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6639_ (.I(_2101_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6640_ (.I(_1047_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6641_ (.A1(_1392_),
    .A2(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6642_ (.A1(_1311_),
    .A2(_1616_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6643_ (.A1(_2102_),
    .A2(_2104_),
    .A3(_2105_),
    .B(_1502_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6644_ (.A1(_1363_),
    .A2(_4130_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6645_ (.I(\as2650.cycle[7] ),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6646_ (.I(_3898_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6647_ (.A1(_2108_),
    .A2(_2109_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6648_ (.A1(_3928_),
    .A2(_3890_),
    .A3(_3929_),
    .A4(_2073_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6649_ (.A1(_2110_),
    .A2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6650_ (.A1(_1038_),
    .A2(_2076_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6651_ (.A1(_1415_),
    .A2(_2112_),
    .A3(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6652_ (.A1(_1059_),
    .A2(_1029_),
    .A3(_1046_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6653_ (.A1(_1633_),
    .A2(_1625_),
    .A3(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6654_ (.A1(_2107_),
    .A2(_2114_),
    .B(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6655_ (.A1(_2088_),
    .A2(_2100_),
    .A3(_2106_),
    .A4(_2117_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6656_ (.I(_2118_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6657_ (.I(_2119_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6658_ (.I(\as2650.addr_buff[0] ),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6659_ (.I(_2121_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6660_ (.I(_2118_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6661_ (.A1(_2122_),
    .A2(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6662_ (.A1(_2071_),
    .A2(_2120_),
    .B(_2124_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6663_ (.I(\as2650.addr_buff[1] ),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6664_ (.I(_2118_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6665_ (.A1(_2125_),
    .A2(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6666_ (.A1(_4225_),
    .A2(_2120_),
    .B(_2127_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6667_ (.I(\as2650.addr_buff[2] ),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6668_ (.A1(_2128_),
    .A2(_2126_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6669_ (.A1(_0308_),
    .A2(_2120_),
    .B(_2129_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6670_ (.I(_1520_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6671_ (.I(\as2650.addr_buff[3] ),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6672_ (.I0(_2130_),
    .I1(_2131_),
    .S(_2119_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6673_ (.I(_2132_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6674_ (.I(_1541_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6675_ (.I(\as2650.addr_buff[4] ),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6676_ (.A1(_2134_),
    .A2(_2126_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6677_ (.A1(_2133_),
    .A2(_2120_),
    .B(_2135_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6678_ (.I(_1535_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6679_ (.I(_3934_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6680_ (.A1(_2137_),
    .A2(_2126_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6681_ (.A1(_2136_),
    .A2(_2123_),
    .B(_2138_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6682_ (.I(_3935_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6683_ (.A1(_2139_),
    .A2(_2119_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6684_ (.A1(_1506_),
    .A2(_2123_),
    .B(_2140_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6685_ (.I(\as2650.addr_buff[7] ),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(_2141_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6687_ (.A1(_2142_),
    .A2(_2119_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6688_ (.A1(_0808_),
    .A2(_2123_),
    .B(_2143_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6689_ (.I(_2074_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6690_ (.A1(_1423_),
    .A2(_2144_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6691_ (.I(_4129_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6692_ (.I(_2146_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6693_ (.A1(_1389_),
    .A2(_1391_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6694_ (.A1(_3941_),
    .A2(_2147_),
    .B(_2148_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6695_ (.A1(_1038_),
    .A2(_1417_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6696_ (.A1(_2149_),
    .A2(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6697_ (.I(_1036_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6698_ (.A1(_1315_),
    .A2(_2152_),
    .A3(_1390_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6699_ (.A1(_3958_),
    .A2(_4056_),
    .A3(_1039_),
    .A4(_1327_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6700_ (.I(_1387_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6701_ (.A1(_1290_),
    .A2(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6702_ (.A1(_1398_),
    .A2(_2153_),
    .A3(_2154_),
    .A4(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6703_ (.A1(_2093_),
    .A2(_2145_),
    .A3(_2151_),
    .A4(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6704_ (.I(_1464_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6705_ (.I(_1672_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6706_ (.A1(_2159_),
    .A2(_2160_),
    .B(_2082_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6707_ (.A1(net24),
    .A2(_2158_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6708_ (.A1(_2158_),
    .A2(_2161_),
    .B(_2162_),
    .C(_1359_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6709_ (.I(_3953_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6710_ (.I(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6711_ (.A1(_2164_),
    .A2(_1410_),
    .A3(_1319_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6712_ (.I(_3955_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6713_ (.I(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6714_ (.I(_2167_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6715_ (.A1(net22),
    .A2(_2165_),
    .B(_2168_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6716_ (.A1(_3870_),
    .A2(_2165_),
    .B(_2169_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6717_ (.I(_1335_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6718_ (.A1(_1031_),
    .A2(_3879_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6719_ (.A1(_2170_),
    .A2(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6720_ (.I(_2172_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6721_ (.I(_2173_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6722_ (.I(_1316_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6723_ (.I(_1470_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6724_ (.I(_1408_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6725_ (.A1(_2175_),
    .A2(_2176_),
    .B(_1290_),
    .C(_2177_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6726_ (.I(_4076_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6727_ (.I(_2179_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6728_ (.A1(_1384_),
    .A2(_3945_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6729_ (.A1(_2180_),
    .A2(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6730_ (.A1(_1026_),
    .A2(_3906_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6731_ (.I(_2183_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6732_ (.A1(_2184_),
    .A2(_1408_),
    .A3(_2153_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6733_ (.A1(_3903_),
    .A2(_1289_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6734_ (.A1(_2183_),
    .A2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6735_ (.A1(_1323_),
    .A2(_2182_),
    .B(_2185_),
    .C(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6736_ (.A1(_2174_),
    .A2(_2178_),
    .B(_2188_),
    .C(_1338_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6737_ (.A1(net23),
    .A2(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6738_ (.I(_2167_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6739_ (.A1(_3882_),
    .A2(_2189_),
    .B(_2190_),
    .C(_2191_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6740_ (.A1(_3991_),
    .A2(_1324_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6741_ (.I(_2192_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6742_ (.I(_2193_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6743_ (.I(_2192_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6744_ (.A1(_4128_),
    .A2(_4136_),
    .A3(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6745_ (.I(_2196_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6746_ (.A1(\as2650.r123[2][0] ),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6747_ (.I(_4154_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6748_ (.A1(_2199_),
    .A2(_1756_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6749_ (.A1(_4127_),
    .A2(_2194_),
    .B(_2198_),
    .C(_2200_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6750_ (.A1(_2199_),
    .A2(_1804_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6751_ (.I(_2196_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6752_ (.A1(\as2650.r123[2][1] ),
    .A2(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6753_ (.A1(_4252_),
    .A2(_2194_),
    .B(_2201_),
    .C(_2203_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6754_ (.A1(_2199_),
    .A2(_1857_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6755_ (.A1(\as2650.r123[2][2] ),
    .A2(_2202_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6756_ (.A1(_0364_),
    .A2(_2194_),
    .B(_2204_),
    .C(_2205_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6757_ (.A1(_2199_),
    .A2(_1895_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6758_ (.A1(\as2650.r123[2][3] ),
    .A2(_2202_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6759_ (.A1(_0457_),
    .A2(_2194_),
    .B(_2206_),
    .C(_2207_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6760_ (.A1(_4155_),
    .A2(_1938_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6761_ (.A1(\as2650.r123[2][4] ),
    .A2(_2202_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6762_ (.A1(_0560_),
    .A2(_2193_),
    .B(_2208_),
    .C(_2209_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6763_ (.A1(_4155_),
    .A2(_1965_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6764_ (.A1(\as2650.r123[2][5] ),
    .A2(_2197_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6765_ (.A1(_0649_),
    .A2(_2193_),
    .B(_2210_),
    .C(_2211_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6766_ (.A1(\as2650.r123[2][6] ),
    .A2(_2197_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6767_ (.A1(_0466_),
    .A2(_1975_),
    .B1(_2193_),
    .B2(_0727_),
    .C(_2212_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6768_ (.A1(_0845_),
    .A2(_2195_),
    .B1(_2197_),
    .B2(\as2650.r123[2][7] ),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6769_ (.A1(_0466_),
    .A2(_1990_),
    .B(_2213_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6770_ (.I(_1044_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6771_ (.I(_1046_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6772_ (.I(_2171_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6773_ (.A1(_1348_),
    .A2(_2214_),
    .A3(_2215_),
    .A4(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6774_ (.A1(_3953_),
    .A2(_1405_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6775_ (.I(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6776_ (.A1(_1400_),
    .A2(_2082_),
    .A3(_2219_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6777_ (.A1(_2217_),
    .A2(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6778_ (.A1(_4048_),
    .A2(_1288_),
    .A3(_1290_),
    .A4(_1393_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6779_ (.A1(_2184_),
    .A2(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6780_ (.A1(_2108_),
    .A2(_3929_),
    .A3(_2073_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6781_ (.A1(_2075_),
    .A2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6782_ (.I(_2225_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6783_ (.A1(_1563_),
    .A2(_2078_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6784_ (.A1(_2226_),
    .A2(_2227_),
    .B(_1463_),
    .C(_2173_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6785_ (.A1(_4134_),
    .A2(_1409_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6786_ (.A1(_1083_),
    .A2(_1309_),
    .A3(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6787_ (.A1(_2031_),
    .A2(_1608_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6788_ (.A1(_1369_),
    .A2(_1380_),
    .B(_1308_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6789_ (.I(_2111_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6790_ (.A1(_1362_),
    .A2(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6791_ (.I(_3930_),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6792_ (.A1(_2108_),
    .A2(_2141_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6793_ (.A1(_1363_),
    .A2(_2235_),
    .A3(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6794_ (.A1(_2231_),
    .A2(_2232_),
    .A3(_2234_),
    .A4(_2237_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6795_ (.A1(_2091_),
    .A2(_2188_),
    .A3(_2230_),
    .A4(_2238_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6796_ (.A1(_2221_),
    .A2(_2223_),
    .A3(_2228_),
    .A4(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6797_ (.A1(_0850_),
    .A2(_1303_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6798_ (.A1(_0635_),
    .A2(_0717_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6799_ (.A1(_3871_),
    .A2(_4070_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6800_ (.A1(_4234_),
    .A2(_0318_),
    .A3(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6801_ (.A1(_0401_),
    .A2(_0547_),
    .A3(_0622_),
    .A4(_2244_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6802_ (.A1(_2242_),
    .A2(_0810_),
    .A3(_2245_),
    .B1(_1302_),
    .B2(_4132_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6803_ (.A1(_2241_),
    .A2(_2246_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6804_ (.A1(_2104_),
    .A2(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6805_ (.I(_1610_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6806_ (.A1(_4048_),
    .A2(_1314_),
    .A3(_2089_),
    .A4(_2113_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6807_ (.A1(_4049_),
    .A2(_2114_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6808_ (.A1(_3932_),
    .A2(_2183_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6809_ (.A1(_3908_),
    .A2(_1404_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6810_ (.A1(_1381_),
    .A2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6811_ (.A1(_1288_),
    .A2(_2183_),
    .A3(_1371_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6812_ (.A1(_2252_),
    .A2(_2254_),
    .B(_2255_),
    .C(_1406_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6813_ (.I(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6814_ (.A1(_3879_),
    .A2(_1054_),
    .A3(_1615_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6815_ (.A1(_0458_),
    .A2(_0853_),
    .B(_2257_),
    .C(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6816_ (.A1(_2250_),
    .A2(_2251_),
    .B(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6817_ (.A1(_2249_),
    .A2(_1618_),
    .B(_2260_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6818_ (.A1(_2240_),
    .A2(_2248_),
    .A3(_2261_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6819_ (.I(_1057_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6820_ (.I(_2263_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6821_ (.A1(_2264_),
    .A2(_2149_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6822_ (.A1(net26),
    .A2(_1349_),
    .A3(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6823_ (.I(_1503_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6824_ (.A1(_3941_),
    .A2(_2149_),
    .B(_2266_),
    .C(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6825_ (.I(_4204_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6826_ (.A1(net26),
    .A2(_2269_),
    .B(_2144_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6827_ (.A1(_1362_),
    .A2(_2074_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6828_ (.I(_2271_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6829_ (.I(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6830_ (.A1(_2096_),
    .A2(_2270_),
    .B(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6831_ (.A1(_2268_),
    .A2(_2274_),
    .B(_2262_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6832_ (.I(_1357_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6833_ (.I(_2276_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6834_ (.A1(net49),
    .A2(_2262_),
    .B(_2275_),
    .C(_2277_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6835_ (.I(net25),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6836_ (.A1(_1054_),
    .A2(_1610_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6837_ (.A1(_1025_),
    .A2(_2279_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6838_ (.A1(_1032_),
    .A2(_3882_),
    .A3(_3960_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6839_ (.A1(_1033_),
    .A2(_2084_),
    .A3(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6840_ (.A1(_2280_),
    .A2(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6841_ (.A1(_2232_),
    .A2(_2283_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6842_ (.A1(_2230_),
    .A2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6843_ (.I(_2037_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6844_ (.A1(_1605_),
    .A2(_2286_),
    .A3(_1294_),
    .B(_2031_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6845_ (.I(_2085_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6846_ (.I(_1332_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6847_ (.A1(_1336_),
    .A2(_3961_),
    .B(_2289_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6848_ (.A1(_2288_),
    .A2(_2290_),
    .B(_2258_),
    .C(_2219_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6849_ (.I(_1633_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6850_ (.A1(_2292_),
    .A2(_1311_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6851_ (.A1(_2083_),
    .A2(_1614_),
    .A3(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6852_ (.A1(_1503_),
    .A2(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6853_ (.A1(_2188_),
    .A2(_2256_),
    .A3(_2291_),
    .A4(_2295_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6854_ (.A1(_2285_),
    .A2(_2287_),
    .A3(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6855_ (.A1(_2248_),
    .A2(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6856_ (.I(_1503_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6857_ (.I(_2083_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6858_ (.A1(net25),
    .A2(_2300_),
    .A3(_2181_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6859_ (.I(_1365_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6860_ (.A1(_2302_),
    .A2(_1296_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6861_ (.I(_2303_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6862_ (.I(_1562_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6863_ (.I(_1611_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6864_ (.A1(net25),
    .A2(_2083_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6865_ (.I(_1034_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6866_ (.I(_2308_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6867_ (.A1(_2309_),
    .A2(_2263_),
    .B(_1042_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6868_ (.A1(_2306_),
    .A2(_2307_),
    .A3(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6869_ (.A1(_2305_),
    .A2(_1612_),
    .B(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6870_ (.A1(_1394_),
    .A2(_2301_),
    .B1(_2304_),
    .B2(_2312_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6871_ (.I(_2313_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6872_ (.A1(_1041_),
    .A2(_2307_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6873_ (.I(_2107_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6874_ (.A1(_2299_),
    .A2(_2314_),
    .B1(_2315_),
    .B2(_2316_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6875_ (.A1(_1609_),
    .A2(_2317_),
    .B(_2298_),
    .C(_2174_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6876_ (.A1(_2278_),
    .A2(_2298_),
    .B(_2318_),
    .C(_2277_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6877_ (.I(_3954_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6878_ (.I(_2272_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6879_ (.A1(_2319_),
    .A2(_3904_),
    .A3(_2079_),
    .A4(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6880_ (.I(_2110_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6881_ (.I(_2322_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6882_ (.A1(_2323_),
    .A2(_2081_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6883_ (.A1(_1463_),
    .A2(_2173_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6884_ (.I(_2075_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6885_ (.A1(_2326_),
    .A2(_2077_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6886_ (.A1(_2325_),
    .A2(_2327_),
    .B(_1434_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6887_ (.A1(_2250_),
    .A2(_2324_),
    .B(_2328_),
    .C(_2092_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6888_ (.A1(_2321_),
    .A2(_2329_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6889_ (.I(_2144_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6890_ (.A1(_2137_),
    .A2(_2331_),
    .B(_2330_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6891_ (.A1(_3976_),
    .A2(_2330_),
    .B(_2332_),
    .C(_2277_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6892_ (.I(_2144_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6893_ (.A1(_2139_),
    .A2(_2333_),
    .B(_2330_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6894_ (.A1(_3975_),
    .A2(_2330_),
    .B(_2334_),
    .C(_2277_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6895_ (.I(_0459_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6896_ (.A1(_4054_),
    .A2(_2146_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6897_ (.A1(_2071_),
    .A2(_2335_),
    .B(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6898_ (.A1(_2289_),
    .A2(_2253_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6899_ (.A1(_2335_),
    .A2(_0444_),
    .A3(_1455_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6900_ (.A1(_3986_),
    .A2(_2252_),
    .A3(_2338_),
    .A4(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6901_ (.A1(_1379_),
    .A2(_1382_),
    .B1(_2254_),
    .B2(_4056_),
    .C(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6902_ (.I(_2341_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6903_ (.I0(_4009_),
    .I1(_2337_),
    .S(_2342_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6904_ (.I(_2343_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6905_ (.I(_1348_),
    .Z(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6906_ (.A1(_1628_),
    .A2(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6907_ (.I(_1482_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6908_ (.A1(_4197_),
    .A2(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6909_ (.A1(_2345_),
    .A2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6910_ (.I0(_4171_),
    .I1(_2348_),
    .S(_2342_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6911_ (.I(_2349_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6912_ (.A1(_0949_),
    .A2(_2147_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6913_ (.A1(_1518_),
    .A2(_1606_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6914_ (.A1(_2350_),
    .A2(_2351_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6915_ (.I(_2341_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6916_ (.I0(_0339_),
    .I1(_2352_),
    .S(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6917_ (.I(_2354_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6918_ (.I(_2335_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6919_ (.I(_2355_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6920_ (.A1(_2130_),
    .A2(_1532_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6921_ (.A1(_1101_),
    .A2(_2356_),
    .B(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6922_ (.I0(_0429_),
    .I1(_2358_),
    .S(_2353_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6923_ (.I(_2359_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6924_ (.I(_1532_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6925_ (.A1(_0519_),
    .A2(_1527_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6926_ (.A1(_2133_),
    .A2(_2360_),
    .B(_2361_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6927_ (.I0(_0485_),
    .I1(_2362_),
    .S(_2353_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6928_ (.I(_2363_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6929_ (.I(_2353_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6930_ (.A1(_2136_),
    .A2(_1482_),
    .B(_1345_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6931_ (.A1(_2364_),
    .A2(_2365_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6932_ (.A1(_0586_),
    .A2(_2364_),
    .B(_2366_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6933_ (.I(_1606_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6934_ (.I0(_1125_),
    .I1(_1506_),
    .S(_2367_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6935_ (.A1(_0683_),
    .A2(_2342_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6936_ (.A1(_2364_),
    .A2(_2368_),
    .B(_2369_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6937_ (.A1(_0808_),
    .A2(_2360_),
    .B(_1526_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6938_ (.A1(_2342_),
    .A2(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6939_ (.A1(_0824_),
    .A2(_2364_),
    .B(_2371_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6940_ (.I(_1357_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6941_ (.I(_2372_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6942_ (.A1(_2373_),
    .A2(_2218_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6943_ (.I(_2163_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6944_ (.I(_2170_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6945_ (.A1(_2375_),
    .A2(_1612_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6946_ (.I(_2101_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6947_ (.A1(_3958_),
    .A2(_3961_),
    .B1(_2377_),
    .B2(_2141_),
    .C(_2263_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6948_ (.A1(_1392_),
    .A2(_2247_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6949_ (.I(_2308_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6950_ (.A1(_2170_),
    .A2(_1383_),
    .A3(_2380_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6951_ (.A1(_2288_),
    .A2(_2379_),
    .A3(_2381_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6952_ (.A1(_2378_),
    .A2(_2382_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6953_ (.I(_2308_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6954_ (.I(_2384_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6955_ (.A1(_1058_),
    .A2(_1479_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6956_ (.A1(_3925_),
    .A2(_1282_),
    .A3(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6957_ (.A1(_1343_),
    .A2(_1305_),
    .B(_2387_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6958_ (.I(_1383_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6959_ (.A1(_2385_),
    .A2(_1390_),
    .B1(_2388_),
    .B2(_2389_),
    .C(_2375_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6960_ (.I(_2179_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6961_ (.I(_2391_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6962_ (.A1(_2105_),
    .A2(_2383_),
    .B1(_2390_),
    .B2(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6963_ (.A1(_2216_),
    .A2(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6964_ (.A1(_2376_),
    .A2(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6965_ (.I(_1562_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6966_ (.I(_2078_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6967_ (.A1(_2396_),
    .A2(_4204_),
    .B(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6968_ (.I(_2380_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6969_ (.A1(_2375_),
    .A2(_2235_),
    .B(_2399_),
    .C(_2346_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6970_ (.I(_1707_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6971_ (.I(_2401_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6972_ (.A1(_2109_),
    .A2(_2269_),
    .B1(_2402_),
    .B2(_2142_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6973_ (.A1(_2154_),
    .A2(_2398_),
    .A3(_2400_),
    .A4(_2403_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6974_ (.A1(_1527_),
    .A2(_1327_),
    .B(_2184_),
    .C(_1504_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6975_ (.A1(_1465_),
    .A2(_2395_),
    .B1(_2404_),
    .B2(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6976_ (.A1(_2374_),
    .A2(_2375_),
    .B1(_1338_),
    .B2(_2406_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6977_ (.A1(_2373_),
    .A2(_2407_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6978_ (.A1(_2374_),
    .A2(_1313_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6979_ (.A1(_2326_),
    .A2(_2224_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6980_ (.I(_2409_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6981_ (.A1(_3907_),
    .A2(_1336_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6982_ (.A1(_2403_),
    .A2(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6983_ (.I(_1040_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6984_ (.A1(_2344_),
    .A2(_2413_),
    .A3(_2398_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6985_ (.A1(_2410_),
    .A2(_2412_),
    .B(_2414_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6986_ (.A1(_2356_),
    .A2(_1327_),
    .B(_2415_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6987_ (.I(_2288_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6988_ (.I(_1617_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6989_ (.A1(_1317_),
    .A2(_2411_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6990_ (.A1(_2418_),
    .A2(_2379_),
    .B1(_2419_),
    .B2(_2413_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6991_ (.I(_1024_),
    .Z(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6992_ (.I(_1614_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6993_ (.A1(_2421_),
    .A2(_2281_),
    .B(_2411_),
    .C(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6994_ (.I(_1312_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6995_ (.A1(_2417_),
    .A2(_2420_),
    .B(_2423_),
    .C(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6996_ (.I(_2391_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6997_ (.A1(_2426_),
    .A2(_2419_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6998_ (.A1(_2355_),
    .A2(_1344_),
    .A3(_2387_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6999_ (.A1(_1344_),
    .A2(_1304_),
    .B(_2427_),
    .C(_2428_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7000_ (.A1(_2267_),
    .A2(_2425_),
    .A3(_2429_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7001_ (.A1(_2159_),
    .A2(_2416_),
    .B(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7002_ (.A1(_2319_),
    .A2(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7003_ (.I(_2276_),
    .Z(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7004_ (.A1(_2408_),
    .A2(_2432_),
    .B(_2433_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7005_ (.I(_2164_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7006_ (.I(_1357_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7007_ (.I(_2385_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7008_ (.I(_2309_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7009_ (.A1(_1037_),
    .A2(_1028_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7010_ (.A1(_1313_),
    .A2(_2170_),
    .B(\as2650.cycle[2] ),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7011_ (.A1(_2437_),
    .A2(_2438_),
    .A3(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7012_ (.A1(_2142_),
    .A2(_2436_),
    .B1(_2281_),
    .B2(_2440_),
    .C(_2264_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7013_ (.A1(_2421_),
    .A2(_1399_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7014_ (.I(_2442_),
    .Z(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7015_ (.I(_2443_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7016_ (.A1(_2300_),
    .A2(_2440_),
    .B(_2444_),
    .C(_2417_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7017_ (.I(_2306_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7018_ (.A1(_3960_),
    .A2(_2073_),
    .A3(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7019_ (.I(_2426_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7020_ (.A1(_2441_),
    .A2(_2445_),
    .B(_2447_),
    .C(_2448_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7021_ (.A1(_3893_),
    .A2(_1028_),
    .B(_2302_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7022_ (.A1(_1366_),
    .A2(_2450_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7023_ (.A1(_1390_),
    .A2(_1416_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7024_ (.A1(_1318_),
    .A2(_2160_),
    .B(_2438_),
    .C(_2439_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7025_ (.A1(_2452_),
    .A2(_2453_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7026_ (.A1(_2451_),
    .A2(_2454_),
    .B(_2273_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7027_ (.A1(_1634_),
    .A2(_2269_),
    .A3(_1410_),
    .A4(_1421_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7028_ (.A1(_2440_),
    .A2(_2456_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7029_ (.I(_2325_),
    .Z(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7030_ (.A1(_2449_),
    .A2(_2455_),
    .B1(_2457_),
    .B2(_2458_),
    .C(_2164_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7031_ (.A1(_2434_),
    .A2(_1037_),
    .B(_2435_),
    .C(_2459_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7032_ (.A1(_3959_),
    .A2(_2438_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7033_ (.I(_2409_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7034_ (.A1(_2109_),
    .A2(_2269_),
    .A3(_2236_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7035_ (.A1(_2461_),
    .A2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7036_ (.I(_2325_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7037_ (.I(_2078_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7038_ (.A1(_2305_),
    .A2(_3984_),
    .B(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7039_ (.A1(_2413_),
    .A2(_2154_),
    .A3(_2464_),
    .A4(_2466_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7040_ (.A1(_2460_),
    .A2(_2463_),
    .B(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7041_ (.A1(_2097_),
    .A2(_2172_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7042_ (.I(_2469_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7043_ (.I(_2470_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7044_ (.I(_2460_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7045_ (.I(_2152_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7046_ (.I(_2473_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7047_ (.A1(_2474_),
    .A2(_2413_),
    .B(_2103_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7048_ (.A1(_1547_),
    .A2(_1322_),
    .A3(_1611_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7049_ (.A1(_1035_),
    .A2(_2103_),
    .B1(_2472_),
    .B2(_2475_),
    .C(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7050_ (.A1(_2471_),
    .A2(_2477_),
    .B(_2374_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7051_ (.I(_1358_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7052_ (.A1(_2434_),
    .A2(_3891_),
    .B1(_2468_),
    .B2(_2478_),
    .C(_2479_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7053_ (.I(\as2650.cycle[4] ),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7054_ (.A1(_2163_),
    .A2(_3891_),
    .A3(_1037_),
    .A4(_1028_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7055_ (.A1(_2480_),
    .A2(_2481_),
    .B(_2168_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7056_ (.A1(_2480_),
    .A2(_2481_),
    .B(_2482_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7057_ (.A1(_2480_),
    .A2(_2481_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7058_ (.A1(\as2650.cycle[5] ),
    .A2(_2483_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7059_ (.A1(_2373_),
    .A2(_2484_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7060_ (.I(_2322_),
    .Z(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7061_ (.I(_2485_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7062_ (.A1(_4140_),
    .A2(_2486_),
    .B1(_2293_),
    .B2(_1349_),
    .C(_2227_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7063_ (.A1(\as2650.cycle[5] ),
    .A2(_2480_),
    .A3(_3959_),
    .A4(_2438_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7064_ (.A1(_2326_),
    .A2(_2488_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7065_ (.A1(_2109_),
    .A2(_2464_),
    .B(_2489_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7066_ (.A1(_2458_),
    .A2(_2487_),
    .B(_2490_),
    .C(_2374_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7067_ (.A1(_2434_),
    .A2(_2326_),
    .B(_2479_),
    .C(_2491_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7068_ (.I(_2402_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7069_ (.I(_2397_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7070_ (.A1(_2356_),
    .A2(_2492_),
    .A3(_2493_),
    .B(_2464_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7071_ (.A1(_2075_),
    .A2(_2488_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7072_ (.A1(_3928_),
    .A2(_2495_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7073_ (.A1(_3885_),
    .A2(_2458_),
    .B1(_2494_),
    .B2(_2496_),
    .C(_2164_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7074_ (.A1(_2434_),
    .A2(_3928_),
    .B(_2479_),
    .C(_2497_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7075_ (.I(_1406_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7076_ (.A1(_1641_),
    .A2(_1352_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7077_ (.A1(\as2650.psu[7] ),
    .A2(_1641_),
    .B(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7078_ (.A1(_2068_),
    .A2(_2498_),
    .B1(_2500_),
    .B2(_1401_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7079_ (.A1(net4),
    .A2(_1401_),
    .A3(_2498_),
    .B(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7080_ (.A1(\as2650.psu[7] ),
    .A2(_2319_),
    .B(_2168_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7081_ (.A1(_2319_),
    .A2(_2502_),
    .B(_2503_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7082_ (.A1(_1362_),
    .A2(_1040_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7083_ (.A1(_1388_),
    .A2(_1391_),
    .B(_2184_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7084_ (.A1(_2223_),
    .A2(_2231_),
    .A3(_2504_),
    .A4(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7085_ (.A1(_2079_),
    .A2(_2476_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7086_ (.A1(_1336_),
    .A2(_3961_),
    .A3(_2086_),
    .B(_2250_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7087_ (.A1(_2220_),
    .A2(_2284_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7088_ (.A1(_2507_),
    .A2(_2508_),
    .A3(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7089_ (.A1(_1035_),
    .A2(_2081_),
    .B(_2103_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7090_ (.A1(_3910_),
    .A2(_1326_),
    .A3(_2241_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7091_ (.I(_2512_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7092_ (.A1(_1036_),
    .A2(_1038_),
    .A3(_1056_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7093_ (.A1(_1035_),
    .A2(_1056_),
    .B1(_2280_),
    .B2(_2514_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7094_ (.A1(_1377_),
    .A2(_2187_),
    .B(_2513_),
    .C(_2515_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7095_ (.A1(_2091_),
    .A2(_2230_),
    .A3(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7096_ (.A1(_1363_),
    .A2(_2511_),
    .B(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7097_ (.A1(_2259_),
    .A2(_2506_),
    .A3(_2510_),
    .A4(_2518_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7098_ (.I(_2519_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7099_ (.I(_2520_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7100_ (.I(_2272_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7101_ (.I(_2522_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7102_ (.I(_1070_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7103_ (.A1(_2180_),
    .A2(_1294_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7104_ (.I(_2525_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7105_ (.I(_2526_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7106_ (.A1(_2179_),
    .A2(_1343_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7107_ (.I(_2528_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7108_ (.I(_0891_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7109_ (.I(_0874_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7110_ (.A1(_0899_),
    .A2(\as2650.stack[1][0] ),
    .B1(\as2650.stack[0][0] ),
    .B2(_2531_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7111_ (.A1(_2530_),
    .A2(_2532_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7112_ (.I(_0875_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7113_ (.I(_1014_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7114_ (.I(_1020_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7115_ (.A1(_2534_),
    .A2(\as2650.stack[3][0] ),
    .B1(\as2650.stack[2][0] ),
    .B2(_2535_),
    .C(_2536_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7116_ (.A1(\as2650.stack[6][0] ),
    .A2(_0906_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7117_ (.A1(_1020_),
    .A2(_2538_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7118_ (.I(_0889_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7119_ (.A1(_2531_),
    .A2(\as2650.stack[5][0] ),
    .B1(\as2650.stack[4][0] ),
    .B2(_0898_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7120_ (.A1(_2540_),
    .A2(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7121_ (.A1(\as2650.stack[7][0] ),
    .A2(_1019_),
    .B(_2539_),
    .C(_2542_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7122_ (.A1(_2533_),
    .A2(_2537_),
    .B(_2543_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7123_ (.I(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7124_ (.I(_2085_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7125_ (.A1(_0459_),
    .A2(_2247_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7126_ (.A1(_2546_),
    .A2(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7127_ (.I(_2548_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7128_ (.A1(_1069_),
    .A2(_2292_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7129_ (.I(_1051_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7130_ (.I(\as2650.addr_buff[0] ),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7131_ (.A1(_4065_),
    .A2(_2551_),
    .B1(_1416_),
    .B2(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7132_ (.A1(_1068_),
    .A2(_4064_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7133_ (.A1(_1030_),
    .A2(_2554_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7134_ (.A1(_1070_),
    .A2(_2443_),
    .B(_2553_),
    .C(_2555_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7135_ (.A1(_1511_),
    .A2(_4004_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7136_ (.A1(net5),
    .A2(_4004_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7137_ (.A1(_2102_),
    .A2(_2558_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7138_ (.A1(_4065_),
    .A2(_2551_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7139_ (.A1(_2557_),
    .A2(_2559_),
    .B(_2560_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7140_ (.A1(_2417_),
    .A2(_2556_),
    .B1(_2561_),
    .B2(_2086_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7141_ (.A1(_2549_),
    .A2(_2550_),
    .B1(_2562_),
    .B2(_2344_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7142_ (.A1(_0459_),
    .A2(_1611_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7143_ (.I(_2564_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7144_ (.A1(_2146_),
    .A2(_1616_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7145_ (.I(_2566_),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7146_ (.A1(_2554_),
    .A2(_2567_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7147_ (.A1(_2524_),
    .A2(_2565_),
    .B(_2568_),
    .C(_2426_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7148_ (.A1(_1636_),
    .A2(_2563_),
    .B(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7149_ (.A1(_2524_),
    .A2(_2527_),
    .B1(_2529_),
    .B2(_2545_),
    .C(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7150_ (.A1(_1383_),
    .A2(_2288_),
    .B(_2379_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7151_ (.I(_2572_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(_2469_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7153_ (.A1(_2573_),
    .A2(_2569_),
    .B(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7154_ (.A1(_2524_),
    .A2(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7155_ (.A1(_2523_),
    .A2(_2571_),
    .B(_2576_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7156_ (.I(_2520_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7157_ (.I(_2167_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7158_ (.A1(_2524_),
    .A2(_2578_),
    .B(_2579_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7159_ (.A1(_2521_),
    .A2(_2577_),
    .B(_2580_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7160_ (.A1(_2259_),
    .A2(_2506_),
    .A3(_2510_),
    .A4(_2518_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7161_ (.I(_2581_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7162_ (.A1(_1082_),
    .A2(_2582_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7163_ (.A1(_1081_),
    .A2(_1069_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7164_ (.A1(_2355_),
    .A2(_2584_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7165_ (.A1(_2215_),
    .A2(_2247_),
    .B(_2585_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7166_ (.I(_1617_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7167_ (.I(_2548_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7168_ (.A1(_1069_),
    .A2(_2292_),
    .B(_1081_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7169_ (.A1(_1081_),
    .A2(_1070_),
    .A3(_1634_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7170_ (.A1(_2587_),
    .A2(_2588_),
    .A3(_2589_),
    .A4(_2590_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7171_ (.I(_2391_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7172_ (.I(_2592_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7173_ (.A1(_2586_),
    .A2(_2591_),
    .B(_2593_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7174_ (.I(_2303_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7175_ (.A1(\as2650.pc[0] ),
    .A2(net5),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7176_ (.A1(_1080_),
    .A2(_1514_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7177_ (.A1(_2596_),
    .A2(_2597_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7178_ (.I(_1051_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7179_ (.I(_2599_),
    .Z(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7180_ (.A1(_4224_),
    .A2(_4085_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7181_ (.A1(_2558_),
    .A2(_2601_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7182_ (.I(_1036_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7183_ (.I(_2603_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7184_ (.A1(_1516_),
    .A2(_2604_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7185_ (.A1(_2600_),
    .A2(_2602_),
    .B(_2605_),
    .C(_1614_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7186_ (.A1(_2125_),
    .A2(_2473_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7187_ (.A1(_1515_),
    .A2(_2309_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7188_ (.A1(_2215_),
    .A2(_2607_),
    .A3(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7189_ (.A1(_2606_),
    .A2(_2609_),
    .B(_1323_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7190_ (.A1(_1633_),
    .A2(_1322_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7191_ (.I(_2611_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7192_ (.A1(_2215_),
    .A2(_2598_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7193_ (.I(_1030_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7194_ (.I(_1615_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7195_ (.I(_2615_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7196_ (.A1(_2612_),
    .A2(_2584_),
    .B1(_2613_),
    .B2(_2614_),
    .C(_2616_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7197_ (.A1(_2587_),
    .A2(_2598_),
    .B1(_2610_),
    .B2(_2617_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7198_ (.A1(_2595_),
    .A2(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7199_ (.I(_2526_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7200_ (.A1(\as2650.stack[7][1] ),
    .A2(_0878_),
    .B(_1019_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7201_ (.I0(\as2650.stack[5][1] ),
    .I1(\as2650.stack[4][1] ),
    .S(_0883_),
    .Z(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7202_ (.A1(\as2650.stack[6][1] ),
    .A2(_2535_),
    .B1(_1015_),
    .B2(_2622_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7203_ (.I(_0872_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7204_ (.I(_0874_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7205_ (.A1(_2624_),
    .A2(\as2650.stack[1][1] ),
    .B1(\as2650.stack[0][1] ),
    .B2(_2625_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7206_ (.A1(_0892_),
    .A2(_2626_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7207_ (.A1(_0903_),
    .A2(\as2650.stack[3][1] ),
    .B1(\as2650.stack[2][1] ),
    .B2(_0906_),
    .C(_2536_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7208_ (.A1(_2621_),
    .A2(_2623_),
    .B1(_2627_),
    .B2(_2628_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7209_ (.I(_2528_),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7210_ (.A1(_2620_),
    .A2(_2584_),
    .B1(_2629_),
    .B2(_2630_),
    .C(_2320_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7211_ (.A1(_2594_),
    .A2(_2619_),
    .A3(_2631_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7212_ (.I(_2520_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7213_ (.A1(_2471_),
    .A2(_2584_),
    .B(_2632_),
    .C(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7214_ (.A1(_2583_),
    .A2(_2634_),
    .B(_2433_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7215_ (.I(_2525_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7216_ (.I(_2635_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7217_ (.A1(_1080_),
    .A2(_1068_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7218_ (.A1(_1092_),
    .A2(_2637_),
    .Z(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7219_ (.I(_2564_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7220_ (.A1(\as2650.pc[1] ),
    .A2(_1512_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7221_ (.A1(\as2650.pc[1] ),
    .A2(_1512_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7222_ (.A1(_2596_),
    .A2(_2640_),
    .B(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7223_ (.A1(\as2650.pc[2] ),
    .A2(net7),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7224_ (.I(_2643_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7225_ (.A1(_2642_),
    .A2(_2644_),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7226_ (.A1(_2421_),
    .A2(_2645_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7227_ (.A1(_2422_),
    .A2(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7228_ (.A1(_2639_),
    .A2(_2638_),
    .B1(_2647_),
    .B2(_2346_),
    .C(_2392_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7229_ (.A1(_1092_),
    .A2(_2589_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7230_ (.A1(_0308_),
    .A2(_2599_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7231_ (.A1(_2128_),
    .A2(_2473_),
    .B(_2650_),
    .C(_1323_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7232_ (.A1(_2421_),
    .A2(_2638_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7233_ (.A1(_2300_),
    .A2(_2646_),
    .A3(_2652_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7234_ (.A1(_1296_),
    .A2(_2546_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7235_ (.A1(_2651_),
    .A2(_2653_),
    .B(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7236_ (.A1(net7),
    .A2(_4216_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7237_ (.A1(_1512_),
    .A2(_4085_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7238_ (.A1(_2558_),
    .A2(_2601_),
    .B(_2657_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7239_ (.A1(_2656_),
    .A2(_2658_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7240_ (.A1(_2656_),
    .A2(_2658_),
    .B(_2102_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7241_ (.A1(_1364_),
    .A2(_1057_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7242_ (.I(_2661_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7243_ (.A1(_1517_),
    .A2(_2603_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7244_ (.A1(_2659_),
    .A2(_2660_),
    .B(_2662_),
    .C(_2663_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7245_ (.A1(_2418_),
    .A2(_2655_),
    .A3(_2664_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7246_ (.A1(_2549_),
    .A2(_2649_),
    .B(_2665_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7247_ (.A1(\as2650.stack[7][2] ),
    .A2(_0878_),
    .B(_1019_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7248_ (.I(_0906_),
    .Z(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7249_ (.I0(\as2650.stack[5][2] ),
    .I1(\as2650.stack[4][2] ),
    .S(_0883_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7250_ (.A1(\as2650.stack[6][2] ),
    .A2(_2668_),
    .B1(_1015_),
    .B2(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7251_ (.A1(_0899_),
    .A2(\as2650.stack[1][2] ),
    .B1(\as2650.stack[0][2] ),
    .B2(_0895_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7252_ (.A1(_0893_),
    .A2(_2671_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7253_ (.A1(_2534_),
    .A2(\as2650.stack[3][2] ),
    .B1(\as2650.stack[2][2] ),
    .B2(_2535_),
    .C(_1021_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7254_ (.A1(_2667_),
    .A2(_2670_),
    .B1(_2672_),
    .B2(_2673_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7255_ (.I(_2186_),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7256_ (.A1(_2648_),
    .A2(_2666_),
    .B1(_2674_),
    .B2(_2675_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7257_ (.A1(_2636_),
    .A2(_2638_),
    .B(_2676_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7258_ (.A1(_2573_),
    .A2(_2648_),
    .B(_2574_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7259_ (.A1(_2638_),
    .A2(_2678_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7260_ (.A1(_2523_),
    .A2(_2677_),
    .B(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7261_ (.A1(_1093_),
    .A2(_2578_),
    .B(_2579_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7262_ (.A1(_2521_),
    .A2(_2680_),
    .B(_2681_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7263_ (.I(_2581_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7264_ (.I(\as2650.pc[3] ),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7265_ (.A1(\as2650.pc[2] ),
    .A2(\as2650.pc[1] ),
    .A3(\as2650.pc[0] ),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7266_ (.A1(_2683_),
    .A2(_2684_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7267_ (.A1(_2683_),
    .A2(net8),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7268_ (.A1(\as2650.pc[3] ),
    .A2(net8),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7269_ (.A1(_2686_),
    .A2(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7270_ (.A1(\as2650.pc[2] ),
    .A2(net7),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7271_ (.I(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7272_ (.A1(_2642_),
    .A2(_2644_),
    .B(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7273_ (.A1(_2688_),
    .A2(_2691_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7274_ (.A1(_2567_),
    .A2(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7275_ (.I(_1312_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7276_ (.A1(_2639_),
    .A2(_2685_),
    .B(_2693_),
    .C(_2694_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7277_ (.I(_2469_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7278_ (.A1(_2573_),
    .A2(_2695_),
    .B(_2696_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7279_ (.I(_2683_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7280_ (.A1(_1068_),
    .A2(_3911_),
    .B(_1092_),
    .C(_1080_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7281_ (.A1(_2698_),
    .A2(_2699_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7282_ (.A1(_1347_),
    .A2(_2263_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7283_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2152_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7284_ (.A1(_0397_),
    .A2(_2101_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7285_ (.A1(_1333_),
    .A2(_2702_),
    .A3(_2703_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7286_ (.A1(_2614_),
    .A2(_2692_),
    .B(_2704_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7287_ (.A1(_2444_),
    .A2(_2685_),
    .B(_2705_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7288_ (.A1(_0304_),
    .A2(_4216_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7289_ (.A1(net8),
    .A2(_0296_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7290_ (.A1(_2707_),
    .A2(_2659_),
    .A3(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7291_ (.A1(_2707_),
    .A2(_2659_),
    .B(_2708_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7292_ (.A1(_2377_),
    .A2(_2710_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7293_ (.A1(_1520_),
    .A2(_2604_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7294_ (.A1(_2709_),
    .A2(_2711_),
    .B(_2712_),
    .C(_2661_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7295_ (.A1(_2701_),
    .A2(_2706_),
    .B(_2713_),
    .C(_2616_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7296_ (.A1(_2549_),
    .A2(_2700_),
    .B(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7297_ (.I(_0898_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7298_ (.A1(_2716_),
    .A2(\as2650.stack[5][3] ),
    .B1(\as2650.stack[4][3] ),
    .B2(_0895_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7299_ (.I(_0890_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7300_ (.A1(\as2650.stack[6][3] ),
    .A2(_2535_),
    .B1(_2718_),
    .B2(\as2650.stack[7][3] ),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7301_ (.A1(_0893_),
    .A2(_2717_),
    .B(_2719_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7302_ (.A1(_0899_),
    .A2(\as2650.stack[1][3] ),
    .B1(\as2650.stack[0][3] ),
    .B2(_0895_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7303_ (.A1(_2534_),
    .A2(\as2650.stack[3][3] ),
    .B1(\as2650.stack[2][3] ),
    .B2(_2540_),
    .C(_2536_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7304_ (.A1(_0893_),
    .A2(_2721_),
    .B(_2722_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7305_ (.A1(_0880_),
    .A2(_2720_),
    .B(_2723_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7306_ (.A1(_2635_),
    .A2(_2685_),
    .B1(_2724_),
    .B2(_2630_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7307_ (.A1(_2695_),
    .A2(_2715_),
    .B(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7308_ (.I(_2470_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7309_ (.A1(_2685_),
    .A2(_2697_),
    .B1(_2726_),
    .B2(_2727_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7310_ (.A1(_2682_),
    .A2(_2728_),
    .B(_2579_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7311_ (.A1(_1100_),
    .A2(_2582_),
    .B(_2729_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7312_ (.I(_1106_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7313_ (.A1(_1347_),
    .A2(_2249_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7314_ (.I(_2731_),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7315_ (.A1(\as2650.pc[4] ),
    .A2(net9),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7316_ (.I(_2733_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7317_ (.A1(_2642_),
    .A2(_2643_),
    .B(_2687_),
    .C(_2690_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7318_ (.A1(_2686_),
    .A2(_2735_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7319_ (.A1(_2734_),
    .A2(_2736_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7320_ (.A1(_1100_),
    .A2(_2684_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7321_ (.A1(_1108_),
    .A2(_2738_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7322_ (.A1(_2732_),
    .A2(_2737_),
    .B1(_2739_),
    .B2(_2565_),
    .C(_2392_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7323_ (.A1(_1100_),
    .A2(_2699_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7324_ (.A1(_1108_),
    .A2(_2741_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7325_ (.A1(_0393_),
    .A2(_0296_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7326_ (.A1(net9),
    .A2(_0406_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7327_ (.A1(_0541_),
    .A2(_0406_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7328_ (.A1(_2743_),
    .A2(_2710_),
    .B(_2744_),
    .C(_2745_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7329_ (.A1(_2744_),
    .A2(_2745_),
    .B(_2743_),
    .C(_2710_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7330_ (.A1(_2377_),
    .A2(_2747_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7331_ (.A1(_1508_),
    .A2(_2551_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7332_ (.A1(_2746_),
    .A2(_2748_),
    .B(_2749_),
    .C(_2661_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7333_ (.A1(\as2650.addr_buff[4] ),
    .A2(_1416_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7334_ (.A1(_4144_),
    .A2(_2737_),
    .B1(_2739_),
    .B2(_2443_),
    .C(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7335_ (.A1(_1509_),
    .A2(_2600_),
    .B(_2752_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7336_ (.A1(_2654_),
    .A2(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7337_ (.A1(_2616_),
    .A2(_2750_),
    .A3(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7338_ (.A1(_2549_),
    .A2(_2742_),
    .B(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7339_ (.I(_2530_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7340_ (.I(_2531_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7341_ (.A1(_2716_),
    .A2(\as2650.stack[1][4] ),
    .B1(\as2650.stack[0][4] ),
    .B2(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7342_ (.A1(_2534_),
    .A2(\as2650.stack[3][4] ),
    .B1(\as2650.stack[2][4] ),
    .B2(_2668_),
    .C(_1021_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7343_ (.A1(_2757_),
    .A2(_2759_),
    .B(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7344_ (.A1(_2716_),
    .A2(\as2650.stack[5][4] ),
    .B1(\as2650.stack[4][4] ),
    .B2(_2758_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7345_ (.A1(\as2650.stack[6][4] ),
    .A2(_2668_),
    .B1(_2718_),
    .B2(\as2650.stack[7][4] ),
    .C(_0880_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7346_ (.A1(_2757_),
    .A2(_2762_),
    .B(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7347_ (.A1(_2761_),
    .A2(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7348_ (.A1(_2526_),
    .A2(_2739_),
    .B1(_2765_),
    .B2(_2630_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7349_ (.A1(_2740_),
    .A2(_2756_),
    .B(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7350_ (.I(_2572_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7351_ (.A1(_2768_),
    .A2(_2740_),
    .B(_2470_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7352_ (.A1(_2574_),
    .A2(_2767_),
    .B1(_2769_),
    .B2(_2739_),
    .C(_2581_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7353_ (.A1(_2730_),
    .A2(_2582_),
    .B(_2770_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7354_ (.A1(_2373_),
    .A2(_2771_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7355_ (.I(_2581_),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7356_ (.A1(_1107_),
    .A2(_1099_),
    .A3(_2684_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7357_ (.A1(_1115_),
    .A2(_2773_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7358_ (.I(_2572_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7359_ (.A1(\as2650.pc[5] ),
    .A2(net1),
    .Z(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7360_ (.A1(_2686_),
    .A2(_2734_),
    .A3(_2735_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7361_ (.A1(_2730_),
    .A2(_0543_),
    .B(_2777_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7362_ (.A1(_2776_),
    .A2(_2778_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7363_ (.A1(_2731_),
    .A2(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7364_ (.I(_2564_),
    .Z(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7365_ (.A1(_2781_),
    .A2(_2774_),
    .B(_1312_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7366_ (.A1(_2775_),
    .A2(_2780_),
    .A3(_2782_),
    .B(_2470_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7367_ (.A1(_2624_),
    .A2(\as2650.stack[1][5] ),
    .B1(\as2650.stack[0][5] ),
    .B2(_2531_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7368_ (.A1(_0892_),
    .A2(_2784_),
    .Z(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7369_ (.A1(_0903_),
    .A2(\as2650.stack[3][5] ),
    .B1(\as2650.stack[2][5] ),
    .B2(_2540_),
    .C(_2536_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7370_ (.A1(_0898_),
    .A2(\as2650.stack[5][5] ),
    .B1(\as2650.stack[4][5] ),
    .B2(_2625_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7371_ (.A1(_0892_),
    .A2(_2787_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7372_ (.A1(\as2650.stack[6][5] ),
    .A2(_2540_),
    .B1(_2718_),
    .B2(\as2650.stack[7][5] ),
    .C(_0880_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7373_ (.A1(_2785_),
    .A2(_2786_),
    .B1(_2788_),
    .B2(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7374_ (.A1(_2730_),
    .A2(_2741_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7375_ (.A1(_1115_),
    .A2(_2791_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7376_ (.A1(_3934_),
    .A2(_1051_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7377_ (.A1(_0616_),
    .A2(_2089_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7378_ (.A1(_1332_),
    .A2(_2793_),
    .A3(_2794_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7379_ (.A1(_2442_),
    .A2(_2774_),
    .B1(_2779_),
    .B2(_4144_),
    .C(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7380_ (.A1(_0615_),
    .A2(_0534_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7381_ (.A1(_2744_),
    .A2(_2746_),
    .A3(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7382_ (.A1(_2744_),
    .A2(_2746_),
    .B(_2797_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7383_ (.A1(_2101_),
    .A2(_2799_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7384_ (.A1(_1535_),
    .A2(_2384_),
    .B1(_2798_),
    .B2(_2800_),
    .C(_2661_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7385_ (.A1(_2701_),
    .A2(_2796_),
    .B(_2801_),
    .C(_2615_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7386_ (.A1(_2548_),
    .A2(_2792_),
    .B(_2802_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7387_ (.A1(_2780_),
    .A2(_2782_),
    .A3(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7388_ (.A1(_2635_),
    .A2(_2774_),
    .B(_2804_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7389_ (.A1(_2675_),
    .A2(_2790_),
    .B(_2805_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7390_ (.A1(_2774_),
    .A2(_2783_),
    .B1(_2806_),
    .B2(_2727_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7391_ (.A1(_2772_),
    .A2(_2807_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7392_ (.I(_2519_),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7393_ (.A1(_1116_),
    .A2(_2809_),
    .B(_2191_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7394_ (.A1(_2808_),
    .A2(_2810_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7395_ (.I(\as2650.pc[6] ),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7396_ (.I(_2811_),
    .Z(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7397_ (.A1(_1115_),
    .A2(_2773_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7398_ (.A1(_2812_),
    .A2(_2813_),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7399_ (.A1(_2624_),
    .A2(\as2650.stack[5][6] ),
    .B1(\as2650.stack[4][6] ),
    .B2(_2625_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7400_ (.A1(\as2650.stack[6][6] ),
    .A2(_1014_),
    .B1(_0890_),
    .B2(\as2650.stack[7][6] ),
    .C(_0879_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7401_ (.A1(_2530_),
    .A2(_2815_),
    .B(_2816_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7402_ (.A1(_2624_),
    .A2(\as2650.stack[1][6] ),
    .B1(\as2650.stack[0][6] ),
    .B2(_2625_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7403_ (.A1(_0903_),
    .A2(\as2650.stack[3][6] ),
    .B1(\as2650.stack[2][6] ),
    .B2(_1014_),
    .C(_1020_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7404_ (.A1(_2530_),
    .A2(_2818_),
    .B(_2819_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7405_ (.A1(_2817_),
    .A2(_2820_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7406_ (.A1(_3885_),
    .A2(_2814_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7407_ (.A1(\as2650.pc[6] ),
    .A2(net2),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7408_ (.I(_2823_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7409_ (.A1(_1114_),
    .A2(net1),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7410_ (.A1(_2777_),
    .A2(_2776_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7411_ (.A1(_1106_),
    .A2(net9),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7412_ (.A1(\as2650.pc[5] ),
    .A2(net1),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7413_ (.A1(_2827_),
    .A2(_2828_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7414_ (.A1(_2825_),
    .A2(_2826_),
    .A3(_2829_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7415_ (.A1(_2824_),
    .A2(_2830_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7416_ (.A1(_1612_),
    .A2(_2831_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7417_ (.A1(_2694_),
    .A2(_2565_),
    .A3(_2832_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7418_ (.I(_4144_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7419_ (.A1(_2834_),
    .A2(_2831_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7420_ (.A1(_2139_),
    .A2(_2604_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7421_ (.A1(_1639_),
    .A2(_2380_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7422_ (.A1(_2836_),
    .A2(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7423_ (.A1(_2175_),
    .A2(_2838_),
    .B(_2701_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7424_ (.A1(_2612_),
    .A2(_2814_),
    .B(_2835_),
    .C(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7425_ (.A1(_1114_),
    .A2(_1106_),
    .A3(_2741_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7426_ (.A1(_2811_),
    .A2(_2841_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7427_ (.A1(_0712_),
    .A2(_0629_),
    .Z(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7428_ (.I(_0615_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7429_ (.A1(_2844_),
    .A2(_0534_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7430_ (.A1(_2845_),
    .A2(_2799_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7431_ (.A1(_2843_),
    .A2(_2846_),
    .Z(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7432_ (.A1(_2600_),
    .A2(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7433_ (.A1(_2843_),
    .A2(_2846_),
    .B(_2848_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7434_ (.I(_2551_),
    .Z(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7435_ (.A1(_1315_),
    .A2(_2546_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7436_ (.I(_2851_),
    .Z(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7437_ (.A1(_1639_),
    .A2(_2850_),
    .B(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7438_ (.I(_2306_),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7439_ (.A1(_2588_),
    .A2(_2842_),
    .B1(_2849_),
    .B2(_2853_),
    .C(_2854_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7440_ (.A1(_2822_),
    .A2(_2833_),
    .B1(_2840_),
    .B2(_2855_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7441_ (.A1(_2636_),
    .A2(_2814_),
    .B1(_2821_),
    .B2(_2529_),
    .C(_2856_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7442_ (.I(_2320_),
    .Z(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7443_ (.A1(_2822_),
    .A2(_2833_),
    .B(_2775_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7444_ (.A1(_2858_),
    .A2(_2859_),
    .B(_2814_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7445_ (.A1(_2523_),
    .A2(_2857_),
    .B(_2860_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7446_ (.A1(_2812_),
    .A2(_2578_),
    .B(_2579_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7447_ (.A1(_2521_),
    .A2(_2861_),
    .B(_2862_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7448_ (.I(\as2650.pc[7] ),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7449_ (.I(_2863_),
    .Z(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7450_ (.A1(_2864_),
    .A2(_2772_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7451_ (.A1(\as2650.pc[6] ),
    .A2(_1114_),
    .A3(_2773_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7452_ (.A1(_2863_),
    .A2(_2866_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7453_ (.A1(_0900_),
    .A2(\as2650.stack[5][7] ),
    .B1(\as2650.stack[4][7] ),
    .B2(_2758_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7454_ (.A1(\as2650.stack[6][7] ),
    .A2(_0907_),
    .B1(_2718_),
    .B2(\as2650.stack[7][7] ),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7455_ (.A1(_2757_),
    .A2(_2868_),
    .B(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7456_ (.A1(_2716_),
    .A2(\as2650.stack[1][7] ),
    .B1(\as2650.stack[0][7] ),
    .B2(_2758_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7457_ (.A1(_0904_),
    .A2(\as2650.stack[3][7] ),
    .B1(\as2650.stack[2][7] ),
    .B2(_2668_),
    .C(_1021_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7458_ (.A1(_2757_),
    .A2(_2871_),
    .B(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7459_ (.A1(_0881_),
    .A2(_2870_),
    .B(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7460_ (.I(_2528_),
    .Z(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7461_ (.A1(_1129_),
    .A2(_1550_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7462_ (.A1(_2811_),
    .A2(_1489_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7463_ (.A1(_2824_),
    .A2(_2830_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7464_ (.A1(_2877_),
    .A2(_2878_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7465_ (.A1(_2876_),
    .A2(_2879_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7466_ (.I(_2384_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7467_ (.A1(_2612_),
    .A2(_2867_),
    .B(_1605_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7468_ (.A1(_2396_),
    .A2(_2881_),
    .B1(_2094_),
    .B2(_2142_),
    .C(_2882_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7469_ (.A1(_2614_),
    .A2(_2880_),
    .B(_2883_),
    .C(_2264_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7470_ (.I(_2548_),
    .Z(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7471_ (.A1(_1123_),
    .A2(_2841_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7472_ (.A1(_1129_),
    .A2(_2886_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7473_ (.A1(_0713_),
    .A2(_0629_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7474_ (.A1(net3),
    .A2(_4103_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7475_ (.A1(_2888_),
    .A2(_2847_),
    .B(_2889_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7476_ (.A1(_2888_),
    .A2(_2847_),
    .A3(_2889_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7477_ (.A1(_2437_),
    .A2(_2890_),
    .A3(_2891_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7478_ (.I(_2599_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7479_ (.A1(_2396_),
    .A2(_2893_),
    .B(_2851_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7480_ (.A1(_2885_),
    .A2(_2887_),
    .B1(_2892_),
    .B2(_2894_),
    .C(_2854_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7481_ (.A1(_2732_),
    .A2(_2880_),
    .B1(_2867_),
    .B2(_2781_),
    .C(_2592_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7482_ (.A1(_2884_),
    .A2(_2895_),
    .B(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7483_ (.A1(_2527_),
    .A2(_2867_),
    .B1(_2874_),
    .B2(_2875_),
    .C(_2897_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7484_ (.A1(_2573_),
    .A2(_2896_),
    .B(_2696_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7485_ (.A1(_2867_),
    .A2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7486_ (.A1(_2523_),
    .A2(_2898_),
    .B(_2900_),
    .C(_2633_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7487_ (.A1(_2865_),
    .A2(_2901_),
    .B(_2433_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7488_ (.A1(_1129_),
    .A2(_2866_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7489_ (.A1(_1158_),
    .A2(_2902_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7490_ (.I(_2903_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7491_ (.I(_2775_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7492_ (.I(_2781_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7493_ (.A1(\as2650.pc[8] ),
    .A2(_0711_),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7494_ (.A1(_2825_),
    .A2(_2829_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7495_ (.A1(_2777_),
    .A2(_2776_),
    .B(_2908_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7496_ (.A1(\as2650.pc[7] ),
    .A2(net2),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7497_ (.A1(_2823_),
    .A2(_2910_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7498_ (.A1(_2863_),
    .A2(_2811_),
    .B(_0712_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7499_ (.A1(_2909_),
    .A2(_2911_),
    .B(_2912_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7500_ (.A1(_2907_),
    .A2(_2913_),
    .Z(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7501_ (.I(_2566_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7502_ (.I(_2302_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7503_ (.A1(_2906_),
    .A2(_2904_),
    .B1(_2914_),
    .B2(_2915_),
    .C(_2916_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7504_ (.A1(_2905_),
    .A2(_2917_),
    .B(_2527_),
    .C(_2273_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7505_ (.A1(_1546_),
    .A2(_4103_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7506_ (.A1(_2919_),
    .A2(_2890_),
    .B(_2603_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7507_ (.A1(_2122_),
    .A2(_2920_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7508_ (.A1(\as2650.pc[8] ),
    .A2(_2863_),
    .A3(_2886_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7509_ (.A1(_2864_),
    .A2(_2886_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7510_ (.A1(_1159_),
    .A2(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7511_ (.A1(_2922_),
    .A2(_2924_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7512_ (.A1(_2122_),
    .A2(_2380_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7513_ (.A1(_2560_),
    .A2(_2926_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7514_ (.A1(_2292_),
    .A2(_2914_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7515_ (.A1(_1634_),
    .A2(_2903_),
    .B(_2928_),
    .C(_2289_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7516_ (.A1(_1317_),
    .A2(_2927_),
    .B(_2929_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7517_ (.I(_2654_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7518_ (.A1(_2588_),
    .A2(_2925_),
    .B1(_2930_),
    .B2(_2931_),
    .C(_2854_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7519_ (.A1(_2852_),
    .A2(_2921_),
    .B(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7520_ (.A1(_0912_),
    .A2(_2529_),
    .B1(_2917_),
    .B2(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7521_ (.I(_2522_),
    .Z(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7522_ (.A1(_2904_),
    .A2(_2918_),
    .B1(_2934_),
    .B2(_2935_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7523_ (.I(_1157_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7524_ (.I(_2166_),
    .Z(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7525_ (.A1(_2937_),
    .A2(_2578_),
    .B(_2938_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7526_ (.A1(_2521_),
    .A2(_2936_),
    .B(_2939_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7527_ (.A1(_2937_),
    .A2(_2902_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7528_ (.A1(_1165_),
    .A2(_2940_),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7529_ (.A1(_1165_),
    .A2(_0712_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7530_ (.A1(_2937_),
    .A2(_0714_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7531_ (.A1(_2907_),
    .A2(_2913_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7532_ (.A1(_2943_),
    .A2(_2944_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7533_ (.A1(_2942_),
    .A2(_2945_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7534_ (.A1(_2906_),
    .A2(_2941_),
    .B1(_2946_),
    .B2(_2915_),
    .C(_2916_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7535_ (.A1(_2905_),
    .A2(_2947_),
    .B(_2858_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7536_ (.A1(_2552_),
    .A2(_2920_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7537_ (.A1(_2125_),
    .A2(_2949_),
    .Z(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7538_ (.A1(_2662_),
    .A2(_2950_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7539_ (.I(\as2650.pc[9] ),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7540_ (.A1(_2952_),
    .A2(_2922_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7541_ (.A1(_2834_),
    .A2(_2946_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7542_ (.I(\as2650.addr_buff[1] ),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7543_ (.A1(_2955_),
    .A2(_2309_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7544_ (.A1(_2605_),
    .A2(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7545_ (.A1(_2444_),
    .A2(_2941_),
    .B1(_2957_),
    .B2(_1317_),
    .C(_2701_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7546_ (.A1(_2588_),
    .A2(_2953_),
    .B1(_2954_),
    .B2(_2958_),
    .C(_2446_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7547_ (.A1(_2951_),
    .A2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7548_ (.A1(_1366_),
    .A2(_2941_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7549_ (.A1(_0927_),
    .A2(_2875_),
    .B1(_2947_),
    .B2(_2960_),
    .C(_2961_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7550_ (.A1(_2941_),
    .A2(_2948_),
    .B1(_2962_),
    .B2(_2935_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7551_ (.A1(_2952_),
    .A2(_2633_),
    .B(_2938_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7552_ (.A1(_2809_),
    .A2(_2963_),
    .B(_2964_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7553_ (.I(\as2650.pc[10] ),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7554_ (.A1(_2965_),
    .A2(_2772_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7555_ (.A1(\as2650.pc[9] ),
    .A2(_1157_),
    .A3(_2902_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7556_ (.A1(_2965_),
    .A2(_2967_),
    .Z(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7557_ (.A1(_2552_),
    .A2(_2955_),
    .A3(_2920_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7558_ (.A1(_2128_),
    .A2(_2969_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7559_ (.A1(_1166_),
    .A2(_2922_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7560_ (.A1(_1172_),
    .A2(_2971_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7561_ (.A1(\as2650.pc[10] ),
    .A2(_1487_),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7562_ (.I(_2973_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7563_ (.A1(_2944_),
    .A2(_2942_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7564_ (.A1(_2952_),
    .A2(_1157_),
    .B(_0713_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7565_ (.A1(_2975_),
    .A2(_2976_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7566_ (.A1(_2974_),
    .A2(_2977_),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7567_ (.A1(\as2650.addr_buff[2] ),
    .A2(_2308_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7568_ (.A1(_2663_),
    .A2(_2979_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7569_ (.A1(_1316_),
    .A2(_2980_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7570_ (.A1(_2611_),
    .A2(_2968_),
    .B(_2981_),
    .C(_2654_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7571_ (.A1(_2834_),
    .A2(_2978_),
    .B(_2982_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7572_ (.A1(_2662_),
    .A2(_2970_),
    .B1(_2972_),
    .B2(_2885_),
    .C(_2983_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7573_ (.A1(_2567_),
    .A2(_2978_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7574_ (.A1(_2565_),
    .A2(_2968_),
    .B(_2985_),
    .C(_2426_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7575_ (.A1(_1636_),
    .A2(_2984_),
    .B(_2986_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7576_ (.A1(_0948_),
    .A2(_2529_),
    .B1(_2968_),
    .B2(_2527_),
    .C(_2987_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7577_ (.A1(_2775_),
    .A2(_2986_),
    .B(_2696_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7578_ (.A1(_2968_),
    .A2(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7579_ (.A1(_2935_),
    .A2(_2988_),
    .B(_2990_),
    .C(_2633_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7580_ (.I(_2276_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7581_ (.A1(_2966_),
    .A2(_2991_),
    .B(_2992_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7582_ (.I(\as2650.pc[11] ),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7583_ (.A1(_1172_),
    .A2(_2967_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7584_ (.A1(_2993_),
    .A2(_2994_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7585_ (.I(_2995_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7586_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7587_ (.A1(_2919_),
    .A2(_2890_),
    .B(_2997_),
    .C(_2152_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7588_ (.A1(_2131_),
    .A2(_2998_),
    .B(_2175_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7589_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2998_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7590_ (.A1(_2389_),
    .A2(_2996_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7591_ (.A1(_2999_),
    .A2(_3000_),
    .B(_3001_),
    .C(_2417_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7592_ (.A1(\as2650.pc[11] ),
    .A2(_1483_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7593_ (.I(_3003_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7594_ (.A1(\as2650.pc[10] ),
    .A2(_1487_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7595_ (.A1(_2974_),
    .A2(_2977_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7596_ (.A1(_3005_),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7597_ (.A1(_3004_),
    .A2(_3007_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7598_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2102_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7599_ (.A1(_2289_),
    .A2(_2712_),
    .A3(_3009_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7600_ (.A1(_2612_),
    .A2(_2995_),
    .B1(_3008_),
    .B2(_2614_),
    .C(_3010_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7601_ (.A1(_1172_),
    .A2(_1165_),
    .A3(_2922_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7602_ (.A1(_1177_),
    .A2(_3012_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7603_ (.A1(_2547_),
    .A2(_3013_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7604_ (.A1(_2379_),
    .A2(_2995_),
    .B(_3014_),
    .C(_2422_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7605_ (.A1(_1532_),
    .A2(_3011_),
    .B(_3015_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7606_ (.A1(_2781_),
    .A2(_2996_),
    .B1(_3008_),
    .B2(_2732_),
    .C(_2592_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7607_ (.I(_3017_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7608_ (.A1(_3002_),
    .A2(_3016_),
    .A3(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7609_ (.A1(_2053_),
    .A2(_2875_),
    .B1(_2996_),
    .B2(_2620_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7610_ (.A1(_3019_),
    .A2(_3020_),
    .B(_2273_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7611_ (.A1(_2858_),
    .A2(_2996_),
    .B(_3021_),
    .C(_2682_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7612_ (.A1(_1178_),
    .A2(_2809_),
    .B(_2191_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7613_ (.A1(_3022_),
    .A2(_3023_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7614_ (.A1(_1185_),
    .A2(_2772_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7615_ (.A1(_2973_),
    .A2(_3004_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7616_ (.A1(_3005_),
    .A2(_2976_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7617_ (.A1(\as2650.pc[11] ),
    .A2(_1488_),
    .B(_3026_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7618_ (.A1(_2975_),
    .A2(_3025_),
    .B(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7619_ (.A1(\as2650.pc[12] ),
    .A2(_0714_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7620_ (.A1(_3028_),
    .A2(_3029_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7621_ (.A1(_2567_),
    .A2(_3030_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7622_ (.A1(_2993_),
    .A2(_2994_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7623_ (.A1(\as2650.pc[12] ),
    .A2(_3032_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7624_ (.A1(_2639_),
    .A2(_3033_),
    .B(_2694_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7625_ (.A1(_3031_),
    .A2(_3034_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7626_ (.A1(_2134_),
    .A2(_3000_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7627_ (.A1(\as2650.pc[12] ),
    .A2(_2993_),
    .A3(_3012_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7628_ (.A1(_1177_),
    .A2(_3012_),
    .B(_1184_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7629_ (.A1(_3037_),
    .A2(_3038_),
    .Z(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7630_ (.A1(\as2650.addr_buff[4] ),
    .A2(_2384_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7631_ (.A1(_2749_),
    .A2(_3040_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7632_ (.A1(_2611_),
    .A2(_3033_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7633_ (.A1(_2834_),
    .A2(_3030_),
    .B1(_3041_),
    .B2(_1607_),
    .C(_3042_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7634_ (.A1(_2885_),
    .A2(_3039_),
    .B1(_3043_),
    .B2(_2931_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7635_ (.A1(_2852_),
    .A2(_3036_),
    .B(_3044_),
    .C(_1636_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _7636_ (.A1(_0973_),
    .A2(_2875_),
    .B1(_3035_),
    .B2(_3045_),
    .C1(_3033_),
    .C2(_2620_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7637_ (.A1(_2768_),
    .A2(_3031_),
    .A3(_3034_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7638_ (.A1(_2858_),
    .A2(_3047_),
    .B(_3033_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7639_ (.A1(_2935_),
    .A2(_3046_),
    .B(_3048_),
    .C(_2520_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7640_ (.A1(_3024_),
    .A2(_3049_),
    .B(_2992_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7641_ (.I(_2893_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7642_ (.A1(_2137_),
    .A2(_3050_),
    .B1(_3000_),
    .B2(_2134_),
    .C(_2852_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7643_ (.A1(_1184_),
    .A2(_1177_),
    .A3(_2994_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7644_ (.A1(_1191_),
    .A2(_3052_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7645_ (.A1(_2137_),
    .A2(_2437_),
    .B1(_2444_),
    .B2(_3053_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7646_ (.A1(\as2650.pc[13] ),
    .A2(_3037_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7647_ (.A1(_1191_),
    .A2(_3037_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7648_ (.A1(_3055_),
    .A2(_3056_),
    .B(_2547_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7649_ (.A1(_2931_),
    .A2(_3054_),
    .B1(_3057_),
    .B2(_2264_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7650_ (.A1(_2768_),
    .A2(_3053_),
    .B(_3058_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7651_ (.A1(_2062_),
    .A2(_2630_),
    .B1(_3053_),
    .B2(_2635_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7652_ (.A1(_2105_),
    .A2(_3051_),
    .A3(_3059_),
    .B(_3060_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7653_ (.A1(_2727_),
    .A2(_2639_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7654_ (.A1(_2471_),
    .A2(_3061_),
    .B1(_3062_),
    .B2(_3053_),
    .C(_2682_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7655_ (.A1(_1191_),
    .A2(_2809_),
    .B(_2168_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7656_ (.A1(_3063_),
    .A2(_3064_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7657_ (.I(\as2650.pc[14] ),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7658_ (.A1(\as2650.pc[13] ),
    .A2(_1184_),
    .A3(_2993_),
    .A4(_2994_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7659_ (.A1(_3065_),
    .A2(_3066_),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7660_ (.A1(\as2650.pc[14] ),
    .A2(_3055_),
    .Z(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7661_ (.A1(_2662_),
    .A2(_2836_),
    .B1(_3068_),
    .B2(_2885_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7662_ (.A1(_2139_),
    .A2(_2385_),
    .B1(_2443_),
    .B2(_3067_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7663_ (.A1(_2422_),
    .A2(_3070_),
    .B(_2931_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7664_ (.A1(_2446_),
    .A2(_3069_),
    .B(_3071_),
    .C(_2424_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7665_ (.A1(_2587_),
    .A2(_2768_),
    .B(_3067_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7666_ (.A1(_2696_),
    .A2(_3072_),
    .B(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7667_ (.A1(_0997_),
    .A2(_2675_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7668_ (.A1(_2471_),
    .A2(_3067_),
    .B1(_3074_),
    .B2(_3075_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7669_ (.A1(_2636_),
    .A2(_3067_),
    .B(_2682_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7670_ (.A1(_3065_),
    .A2(_2582_),
    .B1(_3076_),
    .B2(_3077_),
    .C(_2479_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7671_ (.I(_2222_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7672_ (.A1(_3870_),
    .A2(_1450_),
    .A3(_4082_),
    .B1(_2279_),
    .B2(_3078_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7673_ (.I(_2097_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7674_ (.A1(_3080_),
    .A2(_1607_),
    .A3(_4049_),
    .A4(_2114_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7675_ (.A1(\as2650.addr_buff[7] ),
    .A2(_3936_),
    .Z(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7676_ (.I(_3082_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7677_ (.A1(_2108_),
    .A2(_3083_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7678_ (.A1(_1502_),
    .A2(_2235_),
    .A3(_3084_),
    .B(_3968_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7679_ (.A1(_1385_),
    .A2(_1322_),
    .A3(_1394_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7680_ (.A1(_1502_),
    .A2(_2235_),
    .B(_3926_),
    .C(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7681_ (.A1(_4049_),
    .A2(_3977_),
    .B(_2225_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7682_ (.A1(_1417_),
    .A2(_3088_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7683_ (.A1(_1421_),
    .A2(_1422_),
    .A3(_1382_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7684_ (.A1(_2090_),
    .A2(_3966_),
    .B(_4137_),
    .C(_1046_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7685_ (.A1(_1083_),
    .A2(_3090_),
    .A3(_3091_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7686_ (.A1(_3089_),
    .A2(_3092_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7687_ (.A1(_2097_),
    .A2(_1039_),
    .B(_2528_),
    .C(_2234_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7688_ (.A1(_1374_),
    .A2(_1412_),
    .A3(_2080_),
    .A4(_2229_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7689_ (.A1(_2092_),
    .A2(_2218_),
    .A3(_3094_),
    .A4(_3095_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7690_ (.A1(_3085_),
    .A2(_3087_),
    .B(_3093_),
    .C(_3096_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7691_ (.A1(_1397_),
    .A2(_3079_),
    .A3(_3081_),
    .A4(_3097_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7692_ (.I(_3098_),
    .Z(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7693_ (.I(_3099_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7694_ (.I(_3098_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7695_ (.I(_1451_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7696_ (.I(_2322_),
    .Z(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7697_ (.A1(_3103_),
    .A2(_4124_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7698_ (.A1(_2402_),
    .A2(_4047_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7699_ (.A1(_2850_),
    .A2(_3104_),
    .A3(_3105_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7700_ (.A1(_3050_),
    .A2(_4037_),
    .B(_3106_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7701_ (.A1(_2344_),
    .A2(_4203_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7702_ (.A1(_3102_),
    .A2(_3107_),
    .B(_3108_),
    .C(_2299_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7703_ (.A1(_0443_),
    .A2(_0523_),
    .A3(_0863_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7704_ (.I(_3110_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7705_ (.A1(_4023_),
    .A2(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7706_ (.A1(_3846_),
    .A2(_1479_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7707_ (.I(_3113_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7708_ (.A1(_0885_),
    .A2(_3114_),
    .B(_2038_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7709_ (.I(_0864_),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7710_ (.A1(_4157_),
    .A2(_2037_),
    .B1(_2544_),
    .B2(_3116_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7711_ (.A1(_3112_),
    .A2(_3115_),
    .B(_3117_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7712_ (.A1(_1530_),
    .A2(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7713_ (.I(_3919_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7714_ (.I(_3120_),
    .Z(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7715_ (.A1(_1531_),
    .A2(_4111_),
    .B(_3119_),
    .C(_3121_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7716_ (.I(_1467_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7717_ (.A1(_3123_),
    .A2(_0291_),
    .B(_1471_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7718_ (.A1(_1622_),
    .A2(_1507_),
    .B1(_3122_),
    .B2(_3124_),
    .C(_2694_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7719_ (.I(_3080_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7720_ (.A1(_2448_),
    .A2(_4070_),
    .B(_3125_),
    .C(_3126_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7721_ (.A1(_3101_),
    .A2(_3109_),
    .A3(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7722_ (.I(_2276_),
    .Z(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7723_ (.A1(_1072_),
    .A2(_3100_),
    .B(_3128_),
    .C(_3129_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7724_ (.I(_3101_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7725_ (.I(_2850_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7726_ (.I(_2107_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7727_ (.I(_2401_),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7728_ (.A1(_3133_),
    .A2(_4245_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7729_ (.A1(_2492_),
    .A2(_4249_),
    .B(_3134_),
    .C(_3131_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7730_ (.A1(_3131_),
    .A2(_4195_),
    .B(_3132_),
    .C(_3135_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7731_ (.I(_1379_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7732_ (.I(_3110_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7733_ (.A1(_0896_),
    .A2(_3138_),
    .B(_0854_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7734_ (.A1(_1443_),
    .A2(_3111_),
    .B(_3139_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7735_ (.A1(_4260_),
    .A2(_2037_),
    .B1(_2629_),
    .B2(_3116_),
    .C(_1494_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7736_ (.A1(_3140_),
    .A2(_3141_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7737_ (.I(_1287_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7738_ (.A1(_1478_),
    .A2(_4202_),
    .B(_3142_),
    .C(_3143_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7739_ (.A1(_3123_),
    .A2(_0392_),
    .B(_3144_),
    .C(_1471_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7740_ (.A1(_1628_),
    .A2(_2176_),
    .B(_3145_),
    .C(_2424_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7741_ (.A1(_2448_),
    .A2(_1763_),
    .B(_3146_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7742_ (.A1(_1472_),
    .A2(_3137_),
    .B1(_3147_),
    .B2(_2159_),
    .C(_3098_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7743_ (.A1(_1086_),
    .A2(_3130_),
    .B1(_3136_),
    .B2(_3148_),
    .C(_2372_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7744_ (.I(_2107_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7745_ (.A1(_3133_),
    .A2(_0331_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7746_ (.A1(_3133_),
    .A2(_0337_),
    .B(_3150_),
    .C(_2474_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7747_ (.A1(_3131_),
    .A2(_0363_),
    .B(_3149_),
    .C(_3151_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7748_ (.I(_3120_),
    .Z(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7749_ (.I(\as2650.overflow ),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7750_ (.I0(_0905_),
    .I1(_3154_),
    .S(_3111_),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7751_ (.I(_0853_),
    .Z(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7752_ (.A1(_0369_),
    .A2(_3156_),
    .B1(_2674_),
    .B2(_0870_),
    .C(_1477_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7753_ (.A1(_2038_),
    .A2(_3155_),
    .B(_3157_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7754_ (.A1(_1495_),
    .A2(_1472_),
    .B(_3158_),
    .C(_3121_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7755_ (.A1(_3153_),
    .A2(_1900_),
    .B(_3159_),
    .C(_1501_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7756_ (.A1(_1519_),
    .A2(_1501_),
    .B(_2155_),
    .C(_3160_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7757_ (.A1(_0318_),
    .A2(_2214_),
    .B1(_1379_),
    .B2(_4223_),
    .C(_3098_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7758_ (.A1(_3152_),
    .A2(_3161_),
    .A3(_3162_),
    .Z(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7759_ (.A1(_1094_),
    .A2(_3100_),
    .B(_3163_),
    .C(_3129_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7760_ (.I(_2437_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7761_ (.A1(_2492_),
    .A2(_0422_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7762_ (.A1(_2323_),
    .A2(_0390_),
    .B(_2436_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7763_ (.I(_1414_),
    .Z(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7764_ (.I(_3167_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7765_ (.A1(_3164_),
    .A2(_0456_),
    .B1(_3165_),
    .B2(_3166_),
    .C(_3168_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7766_ (.I0(_1554_),
    .I1(_4016_),
    .S(_3110_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7767_ (.A1(_0472_),
    .A2(_3156_),
    .B(_4207_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7768_ (.A1(_3116_),
    .A2(_2724_),
    .B1(_3170_),
    .B2(_2038_),
    .C(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7769_ (.A1(_1530_),
    .A2(_4223_),
    .B(_3172_),
    .C(_3120_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7770_ (.A1(_3121_),
    .A2(_0614_),
    .B(_3173_),
    .C(_1411_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7771_ (.A1(_2130_),
    .A2(_1501_),
    .B(_2155_),
    .C(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7772_ (.A1(_0401_),
    .A2(_1625_),
    .B1(_1423_),
    .B2(_1900_),
    .C(_3175_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7773_ (.A1(_3101_),
    .A2(_3169_),
    .A3(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7774_ (.A1(_1101_),
    .A2(_3100_),
    .B(_3177_),
    .C(_3129_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7775_ (.A1(_2486_),
    .A2(_0518_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7776_ (.A1(_2492_),
    .A2(_0557_),
    .B(_3050_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7777_ (.A1(_3164_),
    .A2(_0511_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7778_ (.A1(_3178_),
    .A2(_3179_),
    .B(_2316_),
    .C(_3180_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7779_ (.A1(_3952_),
    .A2(_3114_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7780_ (.A1(\as2650.psu[4] ),
    .A2(_3111_),
    .B(_3116_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7781_ (.A1(_0865_),
    .A2(_2765_),
    .B1(_3182_),
    .B2(_3183_),
    .C(_2286_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7782_ (.A1(_1186_),
    .A2(_2286_),
    .B(_3184_),
    .C(_1495_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7783_ (.A1(_1531_),
    .A2(_1900_),
    .B(_3185_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7784_ (.A1(_3153_),
    .A2(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7785_ (.A1(_3123_),
    .A2(_1474_),
    .B(_1408_),
    .C(_2176_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7786_ (.I(_1509_),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7787_ (.A1(_1473_),
    .A2(_1423_),
    .B1(_1389_),
    .B2(_3189_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7788_ (.A1(_0547_),
    .A2(_2214_),
    .B1(_3187_),
    .B2(_3188_),
    .C(_3190_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7789_ (.A1(_3181_),
    .A2(_3191_),
    .B(_3099_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7790_ (.A1(_1109_),
    .A2(_3130_),
    .B(_3192_),
    .C(_3129_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7791_ (.A1(_3103_),
    .A2(_0643_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7792_ (.A1(_2323_),
    .A2(_1940_),
    .B(_3193_),
    .C(_2399_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7793_ (.A1(_3164_),
    .A2(_0611_),
    .B(_3168_),
    .C(_3194_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7794_ (.A1(_1464_),
    .A2(_0622_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7795_ (.A1(_3143_),
    .A2(_0805_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7796_ (.A1(\as2650.psu[5] ),
    .A2(_3138_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7797_ (.A1(\as2650.psl[5] ),
    .A2(_3113_),
    .B(_0855_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7798_ (.A1(_0528_),
    .A2(_3156_),
    .B1(_2790_),
    .B2(_0851_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7799_ (.A1(_3198_),
    .A2(_3199_),
    .B(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7800_ (.I0(_0413_),
    .I1(_3201_),
    .S(_1494_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7801_ (.A1(_3121_),
    .A2(_3202_),
    .B(_1471_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7802_ (.A1(_2136_),
    .A2(_1507_),
    .B1(_3197_),
    .B2(_3203_),
    .C(_2392_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7803_ (.A1(_2177_),
    .A2(_3196_),
    .B(_3204_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7804_ (.A1(_0540_),
    .A2(_3137_),
    .B(_3195_),
    .C(_3205_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7805_ (.A1(_3099_),
    .A2(_3206_),
    .B(_2938_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7806_ (.A1(_1117_),
    .A2(_3100_),
    .B(_3207_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7807_ (.A1(_3164_),
    .A2(_1976_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7808_ (.A1(_2323_),
    .A2(_0706_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7809_ (.A1(_2486_),
    .A2(_0709_),
    .B(_3209_),
    .C(_3050_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7810_ (.A1(_3132_),
    .A2(_3208_),
    .A3(_3210_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7811_ (.I(net27),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7812_ (.A1(_1361_),
    .A2(_3110_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7813_ (.A1(_3212_),
    .A2(_3138_),
    .B(_3213_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7814_ (.A1(_1197_),
    .A2(_3156_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7815_ (.A1(_0864_),
    .A2(_2821_),
    .B(_3215_),
    .C(_1493_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7816_ (.A1(_0855_),
    .A2(_3214_),
    .B(_3216_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7817_ (.A1(_1477_),
    .A2(_0540_),
    .B(_3217_),
    .C(_1467_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7818_ (.A1(_3143_),
    .A2(_4110_),
    .B(_3218_),
    .C(_1470_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7819_ (.A1(_1485_),
    .A2(_1507_),
    .B(_3219_),
    .C(_2592_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7820_ (.A1(_2593_),
    .A2(_2242_),
    .B(_3220_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7821_ (.A1(_0690_),
    .A2(_3137_),
    .B1(_3221_),
    .B2(_2267_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7822_ (.A1(_3211_),
    .A2(_3222_),
    .B(_3099_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7823_ (.I(_1358_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7824_ (.A1(_1125_),
    .A2(_3130_),
    .B(_3223_),
    .C(_3224_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7825_ (.A1(_3133_),
    .A2(_0822_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7826_ (.A1(_2486_),
    .A2(_0803_),
    .B(_2474_),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7827_ (.A1(_3131_),
    .A2(_0844_),
    .B1(_3225_),
    .B2(_3226_),
    .C(_3149_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7828_ (.A1(_0810_),
    .A2(_1625_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7829_ (.A1(\as2650.psu[7] ),
    .A2(_3114_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7830_ (.A1(_1299_),
    .A2(_3114_),
    .B(_3229_),
    .C(_0856_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7831_ (.A1(_1957_),
    .A2(_2286_),
    .B(_1494_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7832_ (.A1(_0870_),
    .A2(_2874_),
    .B(_3231_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7833_ (.A1(_3230_),
    .A2(_3232_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7834_ (.A1(_1497_),
    .A2(_3233_),
    .B(_1469_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7835_ (.A1(_1641_),
    .A2(_2176_),
    .B(_2177_),
    .C(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7836_ (.A1(_1457_),
    .A2(_3137_),
    .B(_3228_),
    .C(_3235_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7837_ (.A1(_3227_),
    .A2(_3236_),
    .B(_3101_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7838_ (.A1(_2068_),
    .A2(_3130_),
    .B(_3237_),
    .C(_3224_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7839_ (.A1(\as2650.stack[6][0] ),
    .A2(_1602_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7840_ (.A1(_1076_),
    .A2(_1600_),
    .B(_3238_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7841_ (.I(_1593_),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7842_ (.A1(\as2650.stack[6][1] ),
    .A2(_1602_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7843_ (.A1(_1089_),
    .A2(_3239_),
    .B(_3240_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7844_ (.I(_1590_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7845_ (.A1(\as2650.stack[6][2] ),
    .A2(_3241_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7846_ (.A1(_1097_),
    .A2(_3239_),
    .B(_3242_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7847_ (.A1(\as2650.stack[6][3] ),
    .A2(_3241_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7848_ (.A1(_1103_),
    .A2(_3239_),
    .B(_3243_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7849_ (.A1(\as2650.stack[6][4] ),
    .A2(_3241_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7850_ (.A1(_1112_),
    .A2(_3239_),
    .B(_3244_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7851_ (.A1(\as2650.stack[6][5] ),
    .A2(_3241_),
    .ZN(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7852_ (.A1(_1120_),
    .A2(_1594_),
    .B(_3245_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7853_ (.A1(\as2650.stack[6][6] ),
    .A2(_1591_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7854_ (.A1(_1127_),
    .A2(_1594_),
    .B(_3246_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7855_ (.A1(\as2650.stack[6][7] ),
    .A2(_1591_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7856_ (.A1(_1131_),
    .A2(_1594_),
    .B(_3247_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7857_ (.I(_1161_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7858_ (.I(_1577_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7859_ (.A1(\as2650.stack[5][8] ),
    .A2(_1586_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7860_ (.A1(_3248_),
    .A2(_3249_),
    .B(_3250_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7861_ (.I(_1168_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7862_ (.I(_1574_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7863_ (.A1(\as2650.stack[5][9] ),
    .A2(_3252_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7864_ (.A1(_3251_),
    .A2(_3249_),
    .B(_3253_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7865_ (.I(_1174_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7866_ (.A1(\as2650.stack[5][10] ),
    .A2(_3252_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7867_ (.A1(_3254_),
    .A2(_3249_),
    .B(_3255_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7868_ (.I(_1181_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7869_ (.A1(\as2650.stack[5][11] ),
    .A2(_3252_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7870_ (.A1(_3256_),
    .A2(_3249_),
    .B(_3257_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7871_ (.I(_1188_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7872_ (.A1(\as2650.stack[5][12] ),
    .A2(_3252_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7873_ (.A1(_3258_),
    .A2(_1578_),
    .B(_3259_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7874_ (.I(_1193_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7875_ (.A1(\as2650.stack[5][13] ),
    .A2(_1575_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7876_ (.A1(_3260_),
    .A2(_1578_),
    .B(_3261_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7877_ (.I(_1199_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7878_ (.A1(\as2650.stack[5][14] ),
    .A2(_1575_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7879_ (.A1(_3262_),
    .A2(_1578_),
    .B(_3263_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7880_ (.I(_1268_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7881_ (.A1(\as2650.stack[4][8] ),
    .A2(_1277_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7882_ (.A1(_3248_),
    .A2(_3264_),
    .B(_3265_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7883_ (.I(_1265_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7884_ (.A1(\as2650.stack[4][9] ),
    .A2(_3266_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7885_ (.A1(_3251_),
    .A2(_3264_),
    .B(_3267_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7886_ (.A1(\as2650.stack[4][10] ),
    .A2(_3266_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7887_ (.A1(_3254_),
    .A2(_3264_),
    .B(_3268_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7888_ (.A1(\as2650.stack[4][11] ),
    .A2(_3266_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7889_ (.A1(_3256_),
    .A2(_3264_),
    .B(_3269_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7890_ (.A1(\as2650.stack[4][12] ),
    .A2(_3266_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7891_ (.A1(_3258_),
    .A2(_1269_),
    .B(_3270_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7892_ (.A1(\as2650.stack[4][13] ),
    .A2(_1266_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7893_ (.A1(_3260_),
    .A2(_1269_),
    .B(_3271_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7894_ (.A1(\as2650.stack[4][14] ),
    .A2(_1266_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7895_ (.A1(_3262_),
    .A2(_1269_),
    .B(_3272_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7896_ (.I(_1251_),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7897_ (.A1(\as2650.stack[3][8] ),
    .A2(_1260_),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7898_ (.A1(_3248_),
    .A2(_3273_),
    .B(_3274_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7899_ (.I(_1248_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7900_ (.A1(\as2650.stack[3][9] ),
    .A2(_3275_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7901_ (.A1(_3251_),
    .A2(_3273_),
    .B(_3276_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7902_ (.A1(\as2650.stack[3][10] ),
    .A2(_3275_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7903_ (.A1(_3254_),
    .A2(_3273_),
    .B(_3277_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7904_ (.A1(\as2650.stack[3][11] ),
    .A2(_3275_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7905_ (.A1(_3256_),
    .A2(_3273_),
    .B(_3278_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7906_ (.A1(\as2650.stack[3][12] ),
    .A2(_3275_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7907_ (.A1(_3258_),
    .A2(_1252_),
    .B(_3279_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7908_ (.A1(\as2650.stack[3][13] ),
    .A2(_1249_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7909_ (.A1(_3260_),
    .A2(_1252_),
    .B(_3280_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7910_ (.A1(\as2650.stack[3][14] ),
    .A2(_1249_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7911_ (.A1(_3262_),
    .A2(_1252_),
    .B(_3281_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7912_ (.A1(_1133_),
    .A2(_1017_),
    .A3(_1264_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7913_ (.I(_3282_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7914_ (.I(_3283_),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7915_ (.I(_3282_),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7916_ (.I(_3285_),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7917_ (.A1(\as2650.stack[7][8] ),
    .A2(_3286_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7918_ (.A1(_3248_),
    .A2(_3284_),
    .B(_3287_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7919_ (.I(_3285_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7920_ (.A1(\as2650.stack[7][9] ),
    .A2(_3288_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7921_ (.A1(_3251_),
    .A2(_3284_),
    .B(_3289_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7922_ (.A1(\as2650.stack[7][10] ),
    .A2(_3288_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7923_ (.A1(_3254_),
    .A2(_3284_),
    .B(_3290_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7924_ (.A1(\as2650.stack[7][11] ),
    .A2(_3288_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7925_ (.A1(_3256_),
    .A2(_3284_),
    .B(_3291_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7926_ (.I(_3283_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7927_ (.A1(\as2650.stack[7][12] ),
    .A2(_3288_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7928_ (.A1(_3258_),
    .A2(_3292_),
    .B(_3293_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7929_ (.I(_3285_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7930_ (.A1(\as2650.stack[7][13] ),
    .A2(_3294_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7931_ (.A1(_3260_),
    .A2(_3292_),
    .B(_3295_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7932_ (.A1(\as2650.stack[7][14] ),
    .A2(_3294_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7933_ (.A1(_3262_),
    .A2(_3292_),
    .B(_3296_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7934_ (.A1(\as2650.stack[7][0] ),
    .A2(_3294_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7935_ (.A1(_1228_),
    .A2(_3292_),
    .B(_3297_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7936_ (.I(_3285_),
    .Z(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7937_ (.A1(\as2650.stack[7][1] ),
    .A2(_3294_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7938_ (.A1(_1232_),
    .A2(_3298_),
    .B(_3299_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7939_ (.I(_3282_),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7940_ (.A1(\as2650.stack[7][2] ),
    .A2(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7941_ (.A1(_1234_),
    .A2(_3298_),
    .B(_3301_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7942_ (.A1(\as2650.stack[7][3] ),
    .A2(_3300_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7943_ (.A1(_1237_),
    .A2(_3298_),
    .B(_3302_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7944_ (.A1(\as2650.stack[7][4] ),
    .A2(_3300_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7945_ (.A1(_1239_),
    .A2(_3298_),
    .B(_3303_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7946_ (.A1(\as2650.stack[7][5] ),
    .A2(_3300_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7947_ (.A1(_1242_),
    .A2(_3286_),
    .B(_3304_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7948_ (.A1(\as2650.stack[7][6] ),
    .A2(_3283_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7949_ (.A1(_1244_),
    .A2(_3286_),
    .B(_3305_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7950_ (.A1(\as2650.stack[7][7] ),
    .A2(_3283_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7951_ (.A1(_1246_),
    .A2(_3286_),
    .B(_3306_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7952_ (.I(net28),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7953_ (.A1(_2248_),
    .A2(_2261_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7954_ (.A1(_1365_),
    .A2(_2603_),
    .A3(_2271_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7955_ (.A1(_3962_),
    .A2(_2086_),
    .B(_2095_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7956_ (.A1(_4140_),
    .A2(_3309_),
    .B1(_3310_),
    .B2(_2216_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7957_ (.A1(_0460_),
    .A2(_2306_),
    .A3(_3311_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7958_ (.A1(_3964_),
    .A2(_2116_),
    .A3(_2187_),
    .A4(_2232_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7959_ (.A1(_2220_),
    .A2(_2230_),
    .A3(_2506_),
    .A4(_3313_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7960_ (.A1(_3308_),
    .A2(_3312_),
    .A3(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7961_ (.I(_3315_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7962_ (.I(_3316_),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7963_ (.A1(_1378_),
    .A2(_2173_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7964_ (.I(_2397_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7965_ (.A1(_3319_),
    .A2(_2554_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7966_ (.I(_2077_),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7967_ (.I(_2112_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7968_ (.I(_3322_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7969_ (.A1(_3977_),
    .A2(_4124_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7970_ (.A1(_2071_),
    .A2(_3324_),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7971_ (.A1(_2141_),
    .A2(_3936_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7972_ (.A1(_4047_),
    .A2(_3326_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7973_ (.A1(_2071_),
    .A2(_3327_),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7974_ (.A1(_3323_),
    .A2(_3325_),
    .B1(_3328_),
    .B2(_2485_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7975_ (.A1(_2233_),
    .A2(_2226_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7976_ (.A1(_3321_),
    .A2(_3329_),
    .B1(_3330_),
    .B2(_3307_),
    .C(_3167_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7977_ (.A1(_2300_),
    .A2(_2615_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7978_ (.A1(_1511_),
    .A2(_2604_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7979_ (.A1(_3307_),
    .A2(_2600_),
    .B(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7980_ (.A1(_2616_),
    .A2(_2554_),
    .B1(_3332_),
    .B2(_3334_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7981_ (.A1(_1333_),
    .A2(_2249_),
    .B(_2303_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7982_ (.I(_3336_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7983_ (.A1(_2304_),
    .A2(_3335_),
    .B1(_3337_),
    .B2(_1071_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7984_ (.A1(_3320_),
    .A2(_3331_),
    .B1(_3338_),
    .B2(_1504_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7985_ (.A1(_1071_),
    .A2(_3318_),
    .B1(_3339_),
    .B2(_2174_),
    .C(_3316_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7986_ (.A1(_3307_),
    .A2(_3317_),
    .B(_3340_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7987_ (.A1(_2433_),
    .A2(_3341_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7988_ (.I(_3315_),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7989_ (.I(_3342_),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7990_ (.I(_3318_),
    .Z(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7991_ (.A1(\as2650.pc[0] ),
    .A2(_4063_),
    .ZN(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7992_ (.A1(_3345_),
    .A2(_2597_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7993_ (.I(_2226_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7994_ (.I(_3322_),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7995_ (.I(_3900_),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7996_ (.I(_3349_),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7997_ (.A1(_4006_),
    .A2(_4166_),
    .A3(_4248_),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7998_ (.A1(_4063_),
    .A2(_4123_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7999_ (.A1(_1556_),
    .A2(_3351_),
    .A3(_3352_),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8000_ (.I(_3349_),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8001_ (.A1(_1516_),
    .A2(_3354_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8002_ (.A1(_3350_),
    .A2(_3353_),
    .B(_3355_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8003_ (.I(_3082_),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8004_ (.A1(_4063_),
    .A2(_4046_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8005_ (.A1(_1556_),
    .A2(_4245_),
    .A3(_3358_),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8006_ (.A1(_1515_),
    .A2(_3357_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8007_ (.A1(_3357_),
    .A2(_3359_),
    .B(_3360_),
    .C(_1708_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8008_ (.A1(_3348_),
    .A2(_3356_),
    .B(_3361_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8009_ (.A1(net53),
    .A2(_3307_),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8010_ (.A1(_2409_),
    .A2(_3363_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8011_ (.A1(_2233_),
    .A2(_2077_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8012_ (.I(_3365_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8013_ (.A1(_3347_),
    .A2(_3362_),
    .B1(_3364_),
    .B2(_3366_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8014_ (.A1(_3319_),
    .A2(_3346_),
    .B(_3367_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8015_ (.I(_2608_),
    .ZN(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8016_ (.A1(_2893_),
    .A2(_3363_),
    .B(_3369_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8017_ (.A1(_2418_),
    .A2(_2598_),
    .B1(_3332_),
    .B2(_3370_),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8018_ (.A1(_1082_),
    .A2(_3337_),
    .B1(_3371_),
    .B2(_2304_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8019_ (.A1(_2316_),
    .A2(_3368_),
    .B1(_3372_),
    .B2(_2299_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8020_ (.I(_2174_),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8021_ (.A1(_1082_),
    .A2(_3344_),
    .B1(_3373_),
    .B2(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8022_ (.A1(net53),
    .A2(_3342_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8023_ (.A1(_3343_),
    .A2(_3375_),
    .B(_3376_),
    .C(_3224_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8024_ (.I(_2145_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8025_ (.I(_3330_),
    .Z(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8026_ (.A1(net53),
    .A2(net28),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8027_ (.A1(net30),
    .A2(_3379_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8028_ (.A1(_3345_),
    .A2(_2640_),
    .B(_2641_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8029_ (.A1(_2644_),
    .A2(_3381_),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8030_ (.I(_3977_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8031_ (.A1(_1513_),
    .A2(_3351_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8032_ (.A1(_1513_),
    .A2(_3351_),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8033_ (.A1(_3352_),
    .A2(_3384_),
    .B(_3385_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8034_ (.A1(_0304_),
    .A2(_0337_),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8035_ (.A1(_3386_),
    .A2(_3387_),
    .B(_3349_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8036_ (.A1(_3386_),
    .A2(_3387_),
    .B(_3388_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8037_ (.A1(_1518_),
    .A2(_3383_),
    .B(_3389_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8038_ (.I(_3326_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8039_ (.A1(_1513_),
    .A2(_4244_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8040_ (.A1(_1514_),
    .A2(_4244_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8041_ (.A1(_3358_),
    .A2(_3392_),
    .B(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8042_ (.A1(_0307_),
    .A2(_0331_),
    .A3(_3394_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8043_ (.A1(_3391_),
    .A2(_3395_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8044_ (.A1(_1518_),
    .A2(_3391_),
    .B(_3396_),
    .C(_2401_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8045_ (.A1(_3348_),
    .A2(_3390_),
    .B(_3397_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8046_ (.A1(_3321_),
    .A2(_3398_),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8047_ (.A1(_3378_),
    .A2(_3380_),
    .B1(_3382_),
    .B2(_3319_),
    .C(_3399_),
    .ZN(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8048_ (.A1(_2893_),
    .A2(_3380_),
    .B(_2650_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8049_ (.A1(_3332_),
    .A2(_3401_),
    .B(_2647_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8050_ (.A1(_1093_),
    .A2(_3337_),
    .B1(_3402_),
    .B2(_2304_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8051_ (.A1(_3168_),
    .A2(_3400_),
    .B1(_3403_),
    .B2(_3126_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8052_ (.A1(_1093_),
    .A2(_3377_),
    .B1(_3404_),
    .B2(_2331_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8053_ (.A1(net30),
    .A2(_3342_),
    .ZN(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8054_ (.A1(_3343_),
    .A2(_3405_),
    .B(_3406_),
    .C(_3224_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8055_ (.I(_3316_),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8056_ (.I(_3407_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8057_ (.I(_3318_),
    .Z(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8058_ (.I(_2409_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8059_ (.A1(_2644_),
    .A2(_3381_),
    .B(_2690_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8060_ (.A1(_2688_),
    .A2(_3411_),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8061_ (.A1(net30),
    .A2(net29),
    .A3(net28),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8062_ (.A1(net31),
    .A2(_3413_),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8063_ (.A1(_0335_),
    .A2(_0336_),
    .B(_0306_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8064_ (.A1(_0305_),
    .A2(_0335_),
    .A3(_0336_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8065_ (.A1(_3386_),
    .A2(_3415_),
    .B(_3416_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8066_ (.A1(_0395_),
    .A2(_0390_),
    .A3(_3417_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8067_ (.A1(_0397_),
    .A2(_3349_),
    .B(_3322_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8068_ (.A1(_3354_),
    .A2(_3418_),
    .B(_3419_),
    .ZN(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8069_ (.A1(_0325_),
    .A2(_0330_),
    .B(_0306_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8070_ (.A1(_0306_),
    .A2(_0325_),
    .A3(_0330_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8071_ (.A1(_3394_),
    .A2(_3421_),
    .B(_3422_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8072_ (.A1(_0395_),
    .A2(_0422_),
    .A3(_3423_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8073_ (.A1(_0397_),
    .A2(_3083_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8074_ (.A1(_3357_),
    .A2(_3424_),
    .B(_3425_),
    .C(_2401_),
    .ZN(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8075_ (.A1(_3420_),
    .A2(_3426_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8076_ (.A1(_3330_),
    .A2(_3414_),
    .B1(_3427_),
    .B2(_2226_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8077_ (.A1(_3410_),
    .A2(_3428_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8078_ (.A1(_3410_),
    .A2(_3412_),
    .B(_3429_),
    .C(_3149_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8079_ (.A1(_2698_),
    .A2(_2389_),
    .A3(_2376_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8080_ (.A1(_2881_),
    .A2(_3414_),
    .B(_2703_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8081_ (.A1(_2175_),
    .A2(_2418_),
    .A3(_3432_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8082_ (.A1(_2214_),
    .A2(_2693_),
    .A3(_3431_),
    .A4(_3433_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8083_ (.A1(_2698_),
    .A2(_2177_),
    .B(_3430_),
    .C(_3434_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8084_ (.A1(_2333_),
    .A2(_3435_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8085_ (.A1(_2698_),
    .A2(_3409_),
    .B(_3436_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8086_ (.A1(net31),
    .A2(_3317_),
    .B(_2938_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8087_ (.A1(_3408_),
    .A2(_3437_),
    .B(_3438_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8088_ (.A1(_2683_),
    .A2(_0393_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8089_ (.A1(_2686_),
    .A2(_3411_),
    .B(_3439_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8090_ (.A1(_2733_),
    .A2(_3440_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8091_ (.A1(_2733_),
    .A2(_3440_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8092_ (.A1(_2465_),
    .A2(_3442_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8093_ (.I(net31),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8094_ (.A1(_3444_),
    .A2(_3413_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8095_ (.A1(net32),
    .A2(_3445_),
    .Z(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8096_ (.A1(_3378_),
    .A2(_3446_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8097_ (.A1(_0394_),
    .A2(_0389_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _8098_ (.A1(_0393_),
    .A2(_0389_),
    .B1(_3386_),
    .B2(_3415_),
    .C(_3416_),
    .ZN(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8099_ (.A1(_3448_),
    .A2(_3449_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8100_ (.A1(_1541_),
    .A2(_0557_),
    .A3(_3450_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8101_ (.A1(_1509_),
    .A2(_3383_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8102_ (.A1(_3383_),
    .A2(_3451_),
    .B(_3452_),
    .C(_3348_),
    .ZN(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8103_ (.I(_3083_),
    .Z(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8104_ (.A1(_0394_),
    .A2(_0421_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _8105_ (.A1(_0394_),
    .A2(_0421_),
    .B1(_3394_),
    .B2(_3421_),
    .C(_3422_),
    .ZN(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8106_ (.A1(_3455_),
    .A2(_3456_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8107_ (.A1(_0543_),
    .A2(_0518_),
    .A3(_3457_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8108_ (.A1(_3454_),
    .A2(_3458_),
    .ZN(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8109_ (.A1(_2133_),
    .A2(_3454_),
    .B(_3459_),
    .C(_2485_),
    .ZN(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8110_ (.A1(_3453_),
    .A2(_3460_),
    .B(_3321_),
    .ZN(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8111_ (.A1(_3441_),
    .A2(_3443_),
    .B(_3447_),
    .C(_3461_),
    .ZN(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8112_ (.A1(_3132_),
    .A2(_3462_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8113_ (.A1(_2377_),
    .A2(_3446_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8114_ (.A1(_2133_),
    .A2(_2881_),
    .B(_3464_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8115_ (.A1(_3332_),
    .A2(_3465_),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8116_ (.A1(_2446_),
    .A2(_2737_),
    .B(_3466_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8117_ (.A1(_1108_),
    .A2(_3337_),
    .B(_3126_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8118_ (.A1(_2916_),
    .A2(_1527_),
    .A3(_3467_),
    .B(_3468_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8119_ (.A1(_3463_),
    .A2(_3469_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8120_ (.A1(_2730_),
    .A2(_3377_),
    .B1(_3470_),
    .B2(_2331_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8121_ (.I(_2166_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8122_ (.A1(net32),
    .A2(_3317_),
    .B(_3472_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8123_ (.A1(_3408_),
    .A2(_3471_),
    .B(_3473_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8124_ (.A1(net32),
    .A2(_3445_),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8125_ (.A1(net52),
    .A2(_3474_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8126_ (.A1(_0541_),
    .A2(_0556_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8127_ (.A1(_0542_),
    .A2(_0556_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8128_ (.A1(_3448_),
    .A2(_3476_),
    .A3(_3449_),
    .B(_3477_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8129_ (.A1(_0617_),
    .A2(_1940_),
    .A3(_3478_),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8130_ (.A1(_0618_),
    .A2(_3354_),
    .B(_3348_),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8131_ (.A1(_3350_),
    .A2(_3479_),
    .B(_3480_),
    .ZN(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8132_ (.A1(_0541_),
    .A2(_0517_),
    .ZN(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8133_ (.A1(_0542_),
    .A2(_0517_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _8134_ (.A1(_3455_),
    .A2(_3482_),
    .A3(_3456_),
    .B(_3483_),
    .ZN(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8135_ (.A1(_0616_),
    .A2(_0643_),
    .A3(_3484_),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8136_ (.A1(_3391_),
    .A2(_3485_),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8137_ (.A1(_2136_),
    .A2(_3391_),
    .B(_3486_),
    .C(_2402_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8138_ (.A1(_3481_),
    .A2(_3487_),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8139_ (.A1(_3378_),
    .A2(_3475_),
    .B1(_3488_),
    .B2(_3347_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8140_ (.A1(_2461_),
    .A2(_3489_),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8141_ (.A1(_2827_),
    .A2(_3442_),
    .ZN(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8142_ (.A1(_2776_),
    .A2(_3491_),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8143_ (.A1(_2493_),
    .A2(_3492_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8144_ (.A1(_3132_),
    .A2(_2333_),
    .A3(_3490_),
    .A4(_3493_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8145_ (.I(_3336_),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8146_ (.A1(_2436_),
    .A2(_3475_),
    .B(_2794_),
    .ZN(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8147_ (.A1(_2389_),
    .A2(_2105_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8148_ (.A1(_1116_),
    .A2(_3495_),
    .B1(_3496_),
    .B2(_3497_),
    .C(_2780_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8149_ (.A1(_2727_),
    .A2(_3498_),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8150_ (.A1(_1116_),
    .A2(_3409_),
    .B(_3494_),
    .C(_3499_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8151_ (.A1(net52),
    .A2(_3317_),
    .B(_3472_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8152_ (.A1(_3408_),
    .A2(_3500_),
    .B(_3501_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8153_ (.I(_3336_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8154_ (.A1(_2160_),
    .A2(_2249_),
    .ZN(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8155_ (.A1(net52),
    .A2(_3474_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8156_ (.A1(net34),
    .A2(_3504_),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8157_ (.A1(_2385_),
    .A2(_3505_),
    .B(_2837_),
    .ZN(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8158_ (.A1(_3503_),
    .A2(_3506_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8159_ (.A1(_2832_),
    .A2(_3507_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8160_ (.A1(_2812_),
    .A2(_3502_),
    .B1(_3508_),
    .B2(_2595_),
    .C(_3126_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8161_ (.A1(_2828_),
    .A2(_3442_),
    .B(_2829_),
    .C(_2825_),
    .ZN(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8162_ (.A1(_2824_),
    .A2(_3510_),
    .Z(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8163_ (.A1(_1487_),
    .A2(_0705_),
    .Z(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8164_ (.A1(_0615_),
    .A2(_0646_),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8165_ (.A1(_2844_),
    .A2(_0646_),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8166_ (.A1(_3478_),
    .A2(_3513_),
    .B(_3514_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8167_ (.A1(_3512_),
    .A2(_3515_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8168_ (.A1(_1489_),
    .A2(_3354_),
    .B(_3322_),
    .ZN(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8169_ (.A1(_3350_),
    .A2(_3516_),
    .B(_3517_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8170_ (.A1(_2844_),
    .A2(_0642_),
    .Z(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8171_ (.A1(_2844_),
    .A2(_0642_),
    .Z(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8172_ (.A1(_3519_),
    .A2(_3484_),
    .B(_3520_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8173_ (.A1(_0714_),
    .A2(_0709_),
    .A3(_3521_),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8174_ (.A1(_1489_),
    .A2(_3083_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8175_ (.A1(_3357_),
    .A2(_3522_),
    .B(_3523_),
    .C(_1708_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8176_ (.A1(_3518_),
    .A2(_3524_),
    .B(_2327_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8177_ (.A1(_3366_),
    .A2(_3505_),
    .B(_3525_),
    .C(_2397_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8178_ (.A1(_3319_),
    .A2(_3511_),
    .B(_3526_),
    .C(_3167_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8179_ (.A1(_3509_),
    .A2(_3527_),
    .B(_2333_),
    .ZN(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8180_ (.A1(_2812_),
    .A2(_3344_),
    .B(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8181_ (.A1(net34),
    .A2(_3342_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8182_ (.A1(_3343_),
    .A2(_3529_),
    .B(_3530_),
    .C(_2435_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8183_ (.A1(_2824_),
    .A2(_3510_),
    .ZN(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8184_ (.A1(_2877_),
    .A2(_3531_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8185_ (.A1(_2876_),
    .A2(_3532_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8186_ (.A1(_1484_),
    .A2(_0706_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8187_ (.A1(_3512_),
    .A2(_3515_),
    .B(_3534_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8188_ (.A1(_1547_),
    .A2(_0822_),
    .A3(_3535_),
    .Z(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8189_ (.A1(_3383_),
    .A2(_3536_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8190_ (.A1(_2305_),
    .A2(_3350_),
    .B(_3323_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8191_ (.A1(_1488_),
    .A2(_0708_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8192_ (.A1(_1488_),
    .A2(_0708_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8193_ (.A1(_3539_),
    .A2(_3521_),
    .B(_3540_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8194_ (.A1(_1547_),
    .A2(_0803_),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8195_ (.A1(_3541_),
    .A2(_3542_),
    .B(_3454_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8196_ (.A1(_3541_),
    .A2(_3542_),
    .B(_3543_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8197_ (.A1(_2396_),
    .A2(_3454_),
    .B(_2485_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8198_ (.A1(_3537_),
    .A2(_3538_),
    .B1(_3544_),
    .B2(_3545_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8199_ (.A1(net34),
    .A2(net33),
    .A3(_3474_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8200_ (.A1(net35),
    .A2(_3547_),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8201_ (.A1(_3366_),
    .A2(_3548_),
    .B(_2465_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8202_ (.A1(_2327_),
    .A2(_3546_),
    .B(_3549_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8203_ (.A1(_2461_),
    .A2(_3533_),
    .B(_3550_),
    .C(_2316_),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8204_ (.A1(_2305_),
    .A2(_2399_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8205_ (.A1(_2399_),
    .A2(_3548_),
    .B(_3552_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8206_ (.A1(_2864_),
    .A2(_3502_),
    .B1(_3497_),
    .B2(_3553_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8207_ (.A1(_2732_),
    .A2(_2880_),
    .B(_3554_),
    .C(_2574_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8208_ (.A1(_2864_),
    .A2(_3344_),
    .B1(_3551_),
    .B2(_3374_),
    .C(_3555_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8209_ (.I(_3316_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8210_ (.A1(net35),
    .A2(_3557_),
    .B(_3472_),
    .ZN(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8211_ (.A1(_3408_),
    .A2(_3556_),
    .B(_3558_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8212_ (.I(_3407_),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8213_ (.I(_3510_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8214_ (.A1(_2911_),
    .A2(_3560_),
    .B(_2912_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8215_ (.A1(_2907_),
    .A2(_3561_),
    .ZN(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8216_ (.I(_3562_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8217_ (.A1(_2907_),
    .A2(_3561_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8218_ (.A1(_2493_),
    .A2(_3563_),
    .A3(_3564_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8219_ (.I(net35),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8220_ (.A1(_3566_),
    .A2(_3547_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8221_ (.A1(net51),
    .A2(_3567_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8222_ (.A1(_0806_),
    .A2(_0802_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8223_ (.A1(_3539_),
    .A2(_3521_),
    .B(_3569_),
    .C(_3540_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8224_ (.A1(_1546_),
    .A2(_0802_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8225_ (.A1(_3082_),
    .A2(_3571_),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8226_ (.A1(_3570_),
    .A2(_3572_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8227_ (.A1(_2552_),
    .A2(_3573_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8228_ (.A1(_0806_),
    .A2(_0821_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8229_ (.A1(_3512_),
    .A2(_3515_),
    .B(_3575_),
    .C(_3534_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8230_ (.A1(_0806_),
    .A2(_0821_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8231_ (.A1(_3900_),
    .A2(_3577_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8232_ (.A1(_3576_),
    .A2(_3578_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8233_ (.A1(_2121_),
    .A2(_3579_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8234_ (.A1(_3103_),
    .A2(_3574_),
    .B1(_3580_),
    .B2(_3323_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8235_ (.A1(_3378_),
    .A2(_3568_),
    .B1(_3581_),
    .B2(_3347_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8236_ (.A1(_2410_),
    .A2(_3582_),
    .B(_3168_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8237_ (.A1(_3565_),
    .A2(_3583_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8238_ (.A1(_2881_),
    .A2(_3568_),
    .B(_3503_),
    .C(_2926_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8239_ (.A1(_2587_),
    .A2(_2914_),
    .B(_3585_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8240_ (.A1(_1159_),
    .A2(_3502_),
    .B1(_3586_),
    .B2(_2595_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8241_ (.A1(_2522_),
    .A2(_3587_),
    .Z(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8242_ (.A1(_2937_),
    .A2(_3344_),
    .B1(_3584_),
    .B2(_3374_),
    .C(_3588_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8243_ (.A1(net51),
    .A2(_3557_),
    .B(_3472_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8244_ (.A1(_3559_),
    .A2(_3589_),
    .B(_3590_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8245_ (.I(_3365_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8246_ (.A1(_3410_),
    .A2(_3591_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8247_ (.A1(net51),
    .A2(_3567_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8248_ (.A1(net37),
    .A2(_3593_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8249_ (.A1(_2121_),
    .A2(_3576_),
    .A3(_3578_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8250_ (.A1(_2955_),
    .A2(_3595_),
    .ZN(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8251_ (.A1(_2121_),
    .A2(_3570_),
    .A3(_3572_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8252_ (.A1(_2955_),
    .A2(_3597_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8253_ (.A1(_3323_),
    .A2(_3596_),
    .B1(_3598_),
    .B2(_3103_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8254_ (.A1(_3347_),
    .A2(_3599_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8255_ (.A1(_3592_),
    .A2(_3594_),
    .B(_3600_),
    .C(_2461_),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8256_ (.I(_2942_),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8257_ (.A1(_2943_),
    .A2(_3602_),
    .A3(_3563_),
    .ZN(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8258_ (.A1(_2943_),
    .A2(_3563_),
    .B(_3602_),
    .ZN(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8259_ (.A1(_2410_),
    .A2(_3604_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8260_ (.A1(_3603_),
    .A2(_3605_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8261_ (.A1(_2367_),
    .A2(_2458_),
    .A3(_3601_),
    .A4(_3606_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8262_ (.A1(_2915_),
    .A2(_2946_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8263_ (.A1(_2474_),
    .A2(_3594_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8264_ (.A1(_2956_),
    .A2(_3609_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8265_ (.A1(_2952_),
    .A2(_3495_),
    .B1(_3497_),
    .B2(_3610_),
    .C(_2522_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8266_ (.A1(_1166_),
    .A2(_3377_),
    .B1(_3608_),
    .B2(_3611_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8267_ (.A1(_3607_),
    .A2(_3612_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8268_ (.I(_2166_),
    .Z(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8269_ (.A1(net37),
    .A2(_3557_),
    .B(_3614_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8270_ (.A1(_3559_),
    .A2(_3613_),
    .B(_3615_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8271_ (.A1(_2122_),
    .A2(_2125_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8272_ (.A1(_3576_),
    .A2(_3578_),
    .B(_1707_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8273_ (.A1(_3570_),
    .A2(_3572_),
    .B(_2322_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8274_ (.A1(_3616_),
    .A2(_3617_),
    .A3(_3618_),
    .ZN(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8275_ (.A1(_2997_),
    .A2(_3617_),
    .A3(_3618_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8276_ (.A1(_3591_),
    .A2(_3620_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8277_ (.A1(_2128_),
    .A2(_3619_),
    .B(_3621_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8278_ (.A1(_1166_),
    .A2(_1159_),
    .B(_1485_),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8279_ (.A1(_3602_),
    .A2(_3563_),
    .ZN(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8280_ (.A1(_3623_),
    .A2(_3624_),
    .B(_2974_),
    .ZN(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8281_ (.A1(_2974_),
    .A2(_3623_),
    .A3(_3624_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8282_ (.A1(_3410_),
    .A2(_3626_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8283_ (.I(net38),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8284_ (.A1(net37),
    .A2(net51),
    .A3(_3567_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8285_ (.A1(_3628_),
    .A2(_3629_),
    .Z(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8286_ (.A1(_3330_),
    .A2(_3630_),
    .Z(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8287_ (.A1(_3625_),
    .A2(_3627_),
    .B(_3167_),
    .C(_3631_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8288_ (.A1(_2473_),
    .A2(_3630_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8289_ (.A1(_2979_),
    .A2(_3633_),
    .ZN(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8290_ (.A1(_2854_),
    .A2(_2978_),
    .B1(_3503_),
    .B2(_3634_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8291_ (.I(_3635_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8292_ (.A1(_2965_),
    .A2(_3495_),
    .B1(_3636_),
    .B2(_2595_),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8293_ (.A1(_3622_),
    .A2(_3632_),
    .B1(_3637_),
    .B2(_1465_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8294_ (.A1(_2965_),
    .A2(_3409_),
    .B1(_3638_),
    .B2(_3374_),
    .ZN(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8295_ (.A1(net38),
    .A2(_3557_),
    .B(_3614_),
    .ZN(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8296_ (.A1(_3559_),
    .A2(_3639_),
    .B(_3640_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8297_ (.A1(_2131_),
    .A2(_3620_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8298_ (.A1(_2997_),
    .A2(_3617_),
    .B(_2233_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8299_ (.A1(_2997_),
    .A2(_3573_),
    .B(_1708_),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8300_ (.A1(_3642_),
    .A2(_3643_),
    .B(_2131_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8301_ (.A1(_3628_),
    .A2(_3629_),
    .ZN(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8302_ (.A1(net39),
    .A2(_3645_),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8303_ (.A1(_3321_),
    .A2(_3644_),
    .B1(_3646_),
    .B2(_3366_),
    .C(_2465_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8304_ (.A1(_3591_),
    .A2(_3641_),
    .B(_3647_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8305_ (.A1(_3005_),
    .A2(_3625_),
    .B(_3003_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8306_ (.I(_3649_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8307_ (.A1(_3005_),
    .A2(_3003_),
    .A3(_3625_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8308_ (.A1(_2493_),
    .A2(_3650_),
    .A3(_3651_),
    .ZN(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8309_ (.A1(_2367_),
    .A2(_2464_),
    .A3(_3648_),
    .A4(_3652_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8310_ (.A1(_2915_),
    .A2(_3008_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8311_ (.A1(_2436_),
    .A2(_3646_),
    .B(_3009_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8312_ (.A1(_1178_),
    .A2(_3495_),
    .B1(_3497_),
    .B2(_3655_),
    .C(_2320_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8313_ (.A1(_3654_),
    .A2(_3656_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8314_ (.A1(_1178_),
    .A2(_3409_),
    .B(_3653_),
    .C(_3657_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8315_ (.A1(net39),
    .A2(_3407_),
    .B(_3614_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8316_ (.A1(_3559_),
    .A2(_3658_),
    .B(_3659_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8317_ (.A1(_2134_),
    .A2(_3641_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8318_ (.A1(_3591_),
    .A2(_3660_),
    .ZN(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8319_ (.A1(net39),
    .A2(_3645_),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8320_ (.A1(net40),
    .A2(_3662_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8321_ (.A1(_3602_),
    .A2(_3025_),
    .A3(_3562_),
    .B(_3027_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8322_ (.A1(_3029_),
    .A2(_3664_),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8323_ (.A1(_3592_),
    .A2(_3663_),
    .B1(_3665_),
    .B2(_2410_),
    .C(_3149_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8324_ (.A1(_2850_),
    .A2(_3663_),
    .ZN(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8325_ (.A1(_2180_),
    .A2(_1316_),
    .A3(_2615_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8326_ (.A1(_3040_),
    .A2(_3667_),
    .B(_3668_),
    .ZN(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8327_ (.A1(_1185_),
    .A2(_3502_),
    .B(_3669_),
    .C(_3031_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8328_ (.I(_3080_),
    .Z(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8329_ (.A1(_3661_),
    .A2(_3666_),
    .B1(_3670_),
    .B2(_3671_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8330_ (.A1(_1185_),
    .A2(_3377_),
    .B1(_3672_),
    .B2(_2331_),
    .ZN(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8331_ (.A1(net40),
    .A2(_3407_),
    .B(_3614_),
    .ZN(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8332_ (.A1(_3343_),
    .A2(_3673_),
    .B(_3674_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8333_ (.A1(_3318_),
    .A2(_2156_),
    .ZN(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8334_ (.A1(_4056_),
    .A2(_2155_),
    .B(_1389_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8335_ (.A1(_4139_),
    .A2(_3964_),
    .A3(_2237_),
    .A4(_3676_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8336_ (.A1(_1463_),
    .A2(_1450_),
    .A3(_2182_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8337_ (.A1(_2092_),
    .A2(_3094_),
    .A3(_3677_),
    .A4(_3678_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8338_ (.A1(_3675_),
    .A2(_2228_),
    .A3(_3679_),
    .ZN(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8339_ (.A1(_3081_),
    .A2(_3680_),
    .ZN(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8340_ (.I(_3681_),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8341_ (.I(_3937_),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8342_ (.I(_3683_),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8343_ (.I(_3683_),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8344_ (.A1(_1072_),
    .A2(_3685_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8345_ (.A1(_3684_),
    .A2(_4203_),
    .B(_3686_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8346_ (.I(_3681_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8347_ (.A1(net41),
    .A2(_3688_),
    .ZN(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8348_ (.A1(_3682_),
    .A2(_3687_),
    .B(_3689_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8349_ (.A1(_1086_),
    .A2(_3685_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8350_ (.A1(_3684_),
    .A2(_1472_),
    .B(_3690_),
    .ZN(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8351_ (.A1(net42),
    .A2(_3688_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8352_ (.A1(_3682_),
    .A2(_3691_),
    .B(_3692_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8353_ (.A1(_1094_),
    .A2(_3685_),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8354_ (.A1(_3684_),
    .A2(_4223_),
    .B(_3693_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8355_ (.A1(net43),
    .A2(_3688_),
    .ZN(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8356_ (.A1(_3682_),
    .A2(_3694_),
    .B(_3695_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8357_ (.A1(_1101_),
    .A2(_3685_),
    .ZN(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8358_ (.A1(_3684_),
    .A2(_0303_),
    .B(_3696_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8359_ (.A1(net44),
    .A2(_3688_),
    .ZN(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8360_ (.A1(_3682_),
    .A2(_3697_),
    .B(_3698_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8361_ (.I(_3681_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8362_ (.I(_3683_),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8363_ (.I(_3683_),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8364_ (.A1(_1109_),
    .A2(_3701_),
    .ZN(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8365_ (.A1(_3700_),
    .A2(_1473_),
    .B(_3702_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8366_ (.I(_3681_),
    .Z(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8367_ (.A1(net45),
    .A2(_3704_),
    .ZN(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8368_ (.A1(_3699_),
    .A2(_3703_),
    .B(_3705_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8369_ (.A1(_1117_),
    .A2(_3701_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8370_ (.A1(_3700_),
    .A2(_1474_),
    .B(_3706_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8371_ (.A1(net19),
    .A2(_3704_),
    .ZN(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8372_ (.A1(_3699_),
    .A2(_3707_),
    .B(_3708_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8373_ (.A1(_1125_),
    .A2(_3701_),
    .ZN(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8374_ (.A1(_3700_),
    .A2(_0805_),
    .B(_3709_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8375_ (.A1(net20),
    .A2(_3704_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8376_ (.A1(_3699_),
    .A2(_3710_),
    .B(_3711_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8377_ (.A1(_2068_),
    .A2(_3701_),
    .ZN(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8378_ (.A1(_3700_),
    .A2(_4110_),
    .B(_3712_),
    .ZN(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8379_ (.A1(net21),
    .A2(_3704_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8380_ (.A1(_3699_),
    .A2(_3713_),
    .B(_3714_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8381_ (.A1(_2130_),
    .A2(_1630_),
    .ZN(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8382_ (.A1(_2916_),
    .A2(_1632_),
    .B(_3715_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8383_ (.A1(_3189_),
    .A2(_1630_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8384_ (.A1(_3671_),
    .A2(_1632_),
    .B(_3716_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8385_ (.I(\as2650.psl[5] ),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8386_ (.A1(_1464_),
    .A2(_1451_),
    .A3(_1318_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8387_ (.A1(_0351_),
    .A2(_2091_),
    .B(_2216_),
    .C(_1388_),
    .ZN(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8388_ (.A1(_1378_),
    .A2(_2229_),
    .A3(_3719_),
    .ZN(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8389_ (.A1(_1333_),
    .A2(_1328_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8390_ (.A1(_3078_),
    .A2(_3721_),
    .B(_1403_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8391_ (.A1(_1375_),
    .A2(_3720_),
    .A3(_3722_),
    .Z(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8392_ (.A1(_2182_),
    .A2(_1417_),
    .A3(_2287_),
    .ZN(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8393_ (.A1(_4097_),
    .A2(_0460_),
    .B1(_3120_),
    .B2(_1530_),
    .C(_2180_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8394_ (.A1(_2147_),
    .A2(_2386_),
    .B(_2498_),
    .C(_3725_),
    .ZN(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8395_ (.A1(_3723_),
    .A2(_3724_),
    .A3(_3726_),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8396_ (.A1(_1346_),
    .A2(_3718_),
    .B(_3727_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8397_ (.A1(_0852_),
    .A2(_1351_),
    .ZN(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8398_ (.I(_3729_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8399_ (.A1(_3730_),
    .A2(_1345_),
    .B(_1478_),
    .ZN(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8400_ (.A1(_1478_),
    .A2(_1473_),
    .B1(_2365_),
    .B2(_3731_),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8401_ (.A1(_3123_),
    .A2(_3732_),
    .B(_3197_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8402_ (.A1(_2299_),
    .A2(_3733_),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8403_ (.A1(_3671_),
    .A2(_0511_),
    .B(_3728_),
    .C(_3734_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8404_ (.A1(_3717_),
    .A2(_3728_),
    .B(_3735_),
    .C(_2435_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8405_ (.A1(_0595_),
    .A2(_1456_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8406_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0595_),
    .B(_3736_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8407_ (.A1(_1428_),
    .A2(_3737_),
    .ZN(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8408_ (.I(_0685_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8409_ (.A1(_3739_),
    .A2(_1976_),
    .ZN(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8410_ (.A1(_0605_),
    .A2(_0610_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8411_ (.A1(_0486_),
    .A2(_0487_),
    .B(_0510_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8412_ (.A1(_0452_),
    .A2(_0455_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8413_ (.A1(_0362_),
    .A2(_0436_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8414_ (.I(_4027_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8415_ (.A1(_3745_),
    .A2(_4036_),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8416_ (.A1(_3745_),
    .A2(_4036_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8417_ (.A1(_4193_),
    .A2(_3747_),
    .B(_4168_),
    .ZN(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8418_ (.A1(_4194_),
    .A2(_3746_),
    .B(_3748_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8419_ (.A1(_0362_),
    .A2(_0436_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8420_ (.A1(_0452_),
    .A2(_0455_),
    .B1(_3744_),
    .B2(_3749_),
    .C(_3750_),
    .ZN(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8421_ (.A1(_0489_),
    .A2(_0509_),
    .ZN(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8422_ (.A1(_3743_),
    .A2(_3751_),
    .B(_3752_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8423_ (.A1(_3741_),
    .A2(_3742_),
    .A3(_3753_),
    .ZN(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8424_ (.A1(_0605_),
    .A2(_0611_),
    .B1(_3739_),
    .B2(_1976_),
    .C(_3754_),
    .ZN(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8425_ (.A1(_1428_),
    .A2(_3737_),
    .B(_2267_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8426_ (.A1(_3738_),
    .A2(_3740_),
    .A3(_3755_),
    .B(_3756_),
    .ZN(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8427_ (.A1(_1622_),
    .A2(_3718_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8428_ (.A1(_3729_),
    .A2(_2336_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8429_ (.A1(_1495_),
    .A2(_2337_),
    .A3(_3759_),
    .ZN(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8430_ (.A1(_1531_),
    .A2(_1457_),
    .B(_3760_),
    .C(_3153_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8431_ (.A1(_3153_),
    .A2(_4203_),
    .B(_3761_),
    .C(_1504_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8432_ (.A1(_3727_),
    .A2(_3758_),
    .A3(_3762_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8433_ (.I(_3763_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8434_ (.A1(_3727_),
    .A2(_3758_),
    .B(_4023_),
    .ZN(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8435_ (.A1(_3757_),
    .A2(_3764_),
    .B(_3765_),
    .C(_2435_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8436_ (.A1(_1451_),
    .A2(_2526_),
    .ZN(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8437_ (.A1(_1519_),
    .A2(_3766_),
    .ZN(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8438_ (.A1(_2514_),
    .A2(_3668_),
    .ZN(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8439_ (.A1(_2272_),
    .A2(_2294_),
    .A3(_2511_),
    .A4(_3768_),
    .ZN(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8440_ (.A1(_2146_),
    .A2(_0444_),
    .A3(_1368_),
    .A4(_0863_),
    .ZN(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8441_ (.A1(_1058_),
    .A2(_3138_),
    .ZN(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8442_ (.A1(_1311_),
    .A2(_1049_),
    .B1(_2546_),
    .B2(_2599_),
    .C(_3771_),
    .ZN(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8443_ (.A1(_2302_),
    .A2(_1605_),
    .B(_3770_),
    .C(_3772_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8444_ (.A1(_2179_),
    .A2(_1318_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8445_ (.A1(_1364_),
    .A2(_2085_),
    .ZN(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8446_ (.A1(_1388_),
    .A2(_1391_),
    .A3(_1616_),
    .A4(_3775_),
    .ZN(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _8447_ (.A1(_3774_),
    .A2(_1339_),
    .A3(_3776_),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8448_ (.A1(_1367_),
    .A2(_3773_),
    .A3(_3777_),
    .ZN(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8449_ (.A1(_2391_),
    .A2(_3143_),
    .A3(_1293_),
    .ZN(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8450_ (.A1(_4135_),
    .A2(_1410_),
    .B1(_2675_),
    .B2(_2335_),
    .C(_2512_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8451_ (.A1(_2287_),
    .A2(_3779_),
    .A3(_3780_),
    .ZN(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8452_ (.A1(_2160_),
    .A2(_1343_),
    .A3(_1329_),
    .A4(_1394_),
    .ZN(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8453_ (.A1(_3769_),
    .A2(_3778_),
    .A3(_3781_),
    .A4(_3782_),
    .ZN(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8454_ (.A1(_3767_),
    .A2(_3783_),
    .ZN(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8455_ (.A1(_1018_),
    .A2(_3784_),
    .ZN(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8456_ (.I(_3783_),
    .Z(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8457_ (.A1(_1352_),
    .A2(_2350_),
    .B(_1295_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8458_ (.A1(_0937_),
    .A2(_1295_),
    .B1(_2352_),
    .B2(_3787_),
    .C(_2593_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8459_ (.A1(_1018_),
    .A2(_0942_),
    .B(_2424_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8460_ (.A1(_1018_),
    .A2(_0942_),
    .B(_3789_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8461_ (.A1(_3788_),
    .A2(_3790_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8462_ (.A1(_3767_),
    .A2(_3786_),
    .A3(_3791_),
    .ZN(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8463_ (.A1(_1359_),
    .A2(_3785_),
    .A3(_3792_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8464_ (.A1(_1628_),
    .A2(_3766_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8465_ (.A1(_3786_),
    .A2(_3793_),
    .B(_0939_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8466_ (.I(_1352_),
    .Z(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8467_ (.A1(_3795_),
    .A2(_2345_),
    .B(_2347_),
    .C(_1344_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8468_ (.A1(_0894_),
    .A2(_1295_),
    .B(_2593_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8469_ (.A1(_2448_),
    .A2(_0894_),
    .B1(_3796_),
    .B2(_3797_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8470_ (.A1(_3786_),
    .A2(_3798_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8471_ (.A1(_3794_),
    .A2(_3799_),
    .B(_2992_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8472_ (.A1(_1622_),
    .A2(_3766_),
    .ZN(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8473_ (.A1(_3786_),
    .A2(_3800_),
    .B(_0943_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8474_ (.A1(_3783_),
    .A2(_3800_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8475_ (.A1(_3795_),
    .A2(_2336_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8476_ (.A1(_2620_),
    .A2(_2337_),
    .A3(_3803_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8477_ (.A1(_0938_),
    .A2(_2636_),
    .B(_3802_),
    .C(_3804_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8478_ (.A1(_2191_),
    .A2(_3801_),
    .A3(_3805_),
    .Z(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8479_ (.I(_3806_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8480_ (.A1(_3080_),
    .A2(_1519_),
    .A3(_2355_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8481_ (.A1(_3774_),
    .A2(_1285_),
    .A3(_3807_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8482_ (.A1(_3723_),
    .A2(_3724_),
    .A3(_3808_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8483_ (.A1(_3730_),
    .A2(_2351_),
    .B(_2350_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8484_ (.A1(_2159_),
    .A2(_3810_),
    .B(_3809_),
    .ZN(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8485_ (.A1(_1428_),
    .A2(_3737_),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8486_ (.A1(_3738_),
    .A2(_3812_),
    .B(_3671_),
    .C(_0830_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8487_ (.A1(_3154_),
    .A2(_3809_),
    .B1(_3811_),
    .B2(_3813_),
    .C(_2372_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8488_ (.A1(_3189_),
    .A2(_2360_),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8489_ (.A1(_2147_),
    .A2(_1370_),
    .ZN(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8490_ (.A1(_2163_),
    .A2(_1607_),
    .A3(_3721_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8491_ (.A1(_1297_),
    .A2(_1348_),
    .B(_2498_),
    .ZN(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8492_ (.A1(_1310_),
    .A2(_3815_),
    .A3(_3816_),
    .A4(_3817_),
    .ZN(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8493_ (.I(_3818_),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8494_ (.A1(_3814_),
    .A2(_3819_),
    .B(_3952_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8495_ (.A1(_3189_),
    .A2(_3102_),
    .A3(_1334_),
    .ZN(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8496_ (.A1(_2361_),
    .A2(_3821_),
    .B(_3819_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8497_ (.I(_3822_),
    .ZN(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8498_ (.A1(_3820_),
    .A2(_3823_),
    .B(_2992_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8499_ (.A1(_2357_),
    .A2(_3819_),
    .B(_4097_),
    .ZN(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8500_ (.A1(_0962_),
    .A2(_2356_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8501_ (.A1(_3730_),
    .A2(_3825_),
    .B(_3819_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8502_ (.A1(_2358_),
    .A2(_3826_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8503_ (.A1(_3824_),
    .A2(_3827_),
    .B(_1360_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8504_ (.A1(_4225_),
    .A2(_3102_),
    .B(_3818_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8505_ (.A1(_3730_),
    .A2(_2347_),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8506_ (.A1(_2348_),
    .A2(_3829_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8507_ (.A1(_1443_),
    .A2(_3828_),
    .B(_2167_),
    .ZN(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8508_ (.A1(_3828_),
    .A2(_3830_),
    .B(_3831_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8509_ (.A1(_1286_),
    .A2(_3771_),
    .B(_2346_),
    .ZN(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8510_ (.A1(_1297_),
    .A2(_0462_),
    .A3(_3816_),
    .A4(_3832_),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8511_ (.A1(_1639_),
    .A2(_2360_),
    .B(_3833_),
    .ZN(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8512_ (.A1(_3102_),
    .A2(_3795_),
    .ZN(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8513_ (.A1(_0998_),
    .A2(_2367_),
    .B1(_3835_),
    .B2(_1506_),
    .ZN(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8514_ (.A1(_3212_),
    .A2(_3834_),
    .B1(_3836_),
    .B2(_3833_),
    .C(_2372_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8515_ (.A1(_1297_),
    .A2(_0462_),
    .A3(_3816_),
    .A4(_3832_),
    .ZN(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8516_ (.A1(_3814_),
    .A2(_3837_),
    .B(\as2650.psu[4] ),
    .ZN(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8517_ (.A1(_3795_),
    .A2(_2361_),
    .ZN(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8518_ (.A1(_2362_),
    .A2(_3833_),
    .A3(_3839_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8519_ (.A1(_3838_),
    .A2(_3840_),
    .B(_1360_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8520_ (.A1(_2357_),
    .A2(_3837_),
    .B(\as2650.psu[3] ),
    .ZN(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8521_ (.A1(_2358_),
    .A2(_3833_),
    .A3(_3835_),
    .ZN(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8522_ (.A1(_3841_),
    .A2(_3842_),
    .B(_1360_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8523_ (.D(_0000_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8524_ (.D(_0001_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8525_ (.D(_0002_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8526_ (.D(_0003_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8527_ (.D(_0004_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8528_ (.D(_0005_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8529_ (.D(_0006_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8530_ (.D(_0007_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8531_ (.D(_0008_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8532_ (.D(_0009_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8533_ (.D(_0010_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8534_ (.D(_0011_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8535_ (.D(_0012_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8536_ (.D(_0013_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8537_ (.D(_0014_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8538_ (.D(_0015_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8539_ (.D(_0016_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8540_ (.D(_0017_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8541_ (.D(_0018_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8542_ (.D(_0019_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8543_ (.D(_0020_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8544_ (.D(_0021_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8545_ (.D(_0022_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8546_ (.D(_0023_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8547_ (.D(_0024_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8548_ (.D(_0025_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8549_ (.D(_0026_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8550_ (.D(_0027_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8551_ (.D(_0028_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8552_ (.D(_0029_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8553_ (.D(_0030_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8554_ (.D(_0031_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8555_ (.D(_0032_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8556_ (.D(_0033_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8557_ (.D(_0034_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8558_ (.D(_0035_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8559_ (.D(_0036_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8560_ (.D(_0037_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8561_ (.D(_0038_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8562_ (.D(_0039_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8563_ (.D(_0040_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8564_ (.D(_0041_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8565_ (.D(_0042_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8566_ (.D(_0043_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8567_ (.D(_0044_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8568_ (.D(_0045_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8569_ (.D(_0046_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8570_ (.D(_0047_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8571_ (.D(_0048_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8572_ (.D(_0049_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8573_ (.D(_0050_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8574_ (.D(_0051_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8575_ (.D(_0052_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8576_ (.D(_0053_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8577_ (.D(_0054_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8578_ (.D(_0055_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8579_ (.D(_0056_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8580_ (.D(_0057_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8581_ (.D(_0058_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8582_ (.D(_0059_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8583_ (.D(_0060_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8584_ (.D(_0061_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8585_ (.D(_0062_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8586_ (.D(_0063_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8587_ (.D(_0064_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8588_ (.D(_0065_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8589_ (.D(_0066_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8590_ (.D(_0067_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8591_ (.D(_0068_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8592_ (.D(_0069_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8593_ (.D(_0070_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8594_ (.D(_0071_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8595_ (.D(_0072_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8596_ (.D(_0073_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8597_ (.D(_0074_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8598_ (.D(_0075_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8599_ (.D(_0076_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8600_ (.D(_0077_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8601_ (.D(_0078_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8602_ (.D(_0079_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8603_ (.D(_0080_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8604_ (.D(_0081_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8605_ (.D(_0082_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8606_ (.D(_0083_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8607_ (.D(_0084_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8608_ (.D(_0085_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8609_ (.D(_0086_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8610_ (.D(_0087_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8611_ (.D(_0088_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8612_ (.D(_0089_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8613_ (.D(_0090_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8614_ (.D(_0091_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8615_ (.D(_0092_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8616_ (.D(_0093_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8617_ (.D(_0094_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8618_ (.D(_0095_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8619_ (.D(_0096_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8620_ (.D(_0097_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8621_ (.D(_0098_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8622_ (.D(_0099_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8623_ (.D(_0100_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8624_ (.D(_0101_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8625_ (.D(_0102_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8626_ (.D(_0103_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8627_ (.D(_0104_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8628_ (.D(_0105_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8629_ (.D(_0106_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8630_ (.D(_0107_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8631_ (.D(_0108_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8632_ (.D(_0109_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8633_ (.D(_0110_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8634_ (.D(_0111_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8635_ (.D(_0112_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8636_ (.D(_0113_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8637_ (.D(_0114_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8638_ (.D(_0115_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8639_ (.D(_0116_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8640_ (.D(_0117_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8641_ (.D(_0118_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8642_ (.D(_0119_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8643_ (.D(_0120_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8644_ (.D(_0121_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8645_ (.D(_0122_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8646_ (.D(_0123_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8647_ (.D(_0124_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8648_ (.D(_0125_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8649_ (.D(_0126_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8650_ (.D(_0127_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8651_ (.D(_0128_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8652_ (.D(_0129_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8653_ (.D(_0130_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8654_ (.D(_0131_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8655_ (.D(_0132_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8656_ (.D(_0133_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8657_ (.D(_0134_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8658_ (.D(_0135_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8659_ (.D(_0136_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8660_ (.D(_0137_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8661_ (.D(_0138_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8662_ (.D(_0139_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8663_ (.D(_0140_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8664_ (.D(_0141_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8665_ (.D(_0142_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8666_ (.D(_0143_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8667_ (.D(_0144_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8668_ (.D(_0145_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8669_ (.D(_0146_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8670_ (.D(_0147_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8671_ (.D(_0148_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8672_ (.D(_0149_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8673_ (.D(_0150_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8674_ (.D(_0151_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8675_ (.D(_0152_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8676_ (.D(_0153_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8677_ (.D(_0154_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8678_ (.D(_0155_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8679_ (.D(_0156_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8680_ (.D(_0157_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8681_ (.D(_0158_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8682_ (.D(_0159_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8683_ (.D(_0160_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8684_ (.D(_0161_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8685_ (.D(_0162_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _8686_ (.D(_0163_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8687_ (.D(_0164_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8688_ (.D(_0165_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8689_ (.D(_0166_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8690_ (.D(_0167_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8691_ (.D(_0168_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8692_ (.D(_0169_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8693_ (.D(_0170_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8694_ (.D(_0171_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8695_ (.D(_0172_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8696_ (.D(_0173_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8697_ (.D(_0174_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8698_ (.D(_0175_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8699_ (.D(_0176_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8700_ (.D(_0177_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8701_ (.D(_0178_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8702_ (.D(_0179_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8703_ (.D(_0180_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8704_ (.D(_0181_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8705_ (.D(_0182_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8706_ (.D(_0183_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8707_ (.D(_0184_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8708_ (.D(_0185_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8709_ (.D(_0186_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8710_ (.D(_0187_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8711_ (.D(_0188_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8712_ (.D(_0189_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8713_ (.D(_0190_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8714_ (.D(_0191_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8715_ (.D(_0192_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8716_ (.D(_0193_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8717_ (.D(_0194_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8718_ (.D(_0195_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8719_ (.D(_0196_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8720_ (.D(_0197_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8721_ (.D(_0198_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8722_ (.D(_0199_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8723_ (.D(_0200_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8724_ (.D(_0201_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8725_ (.D(_0202_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8726_ (.D(_0203_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8727_ (.D(_0204_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8728_ (.D(_0205_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8729_ (.D(_0206_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8730_ (.D(_0207_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8731_ (.D(_0208_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8732_ (.D(_0209_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8733_ (.D(_0210_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8734_ (.D(_0211_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8735_ (.D(_0212_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8736_ (.D(_0213_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8737_ (.D(_0214_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8738_ (.D(_0215_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8739_ (.D(_0216_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8740_ (.D(_0217_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8741_ (.D(_0218_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8742_ (.D(_0219_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8743_ (.D(_0220_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8744_ (.D(_0221_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8745_ (.D(_0222_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8746_ (.D(_0223_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8747_ (.D(_0224_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8748_ (.D(_0225_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8749_ (.D(_0226_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8750_ (.D(_0227_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8751_ (.D(_0228_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8752_ (.D(_0229_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8753_ (.D(_0230_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8754_ (.D(_0231_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8755_ (.D(_0232_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8756_ (.D(_0233_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8757_ (.D(_0234_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8758_ (.D(_0235_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8759_ (.D(_0236_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8760_ (.D(_0237_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8761_ (.D(_0238_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8762_ (.D(_0239_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8763_ (.D(_0240_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8764_ (.D(_0241_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8765_ (.D(_0242_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8766_ (.D(_0243_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8767_ (.D(_0244_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8768_ (.D(_0245_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8769_ (.D(_0246_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8770_ (.D(_0247_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8771_ (.D(_0248_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8772_ (.D(_0249_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8773_ (.D(_0250_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8774_ (.D(_0251_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8775_ (.D(_0252_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8776_ (.D(_0253_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8777_ (.D(_0254_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8778_ (.D(_0255_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8779_ (.D(_0256_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8780_ (.D(_0257_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8781_ (.D(_0258_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8782_ (.D(_0259_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8783_ (.D(_0260_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8784_ (.D(_0261_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8785_ (.D(_0262_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8786_ (.D(_0263_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8787_ (.D(_0264_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8788_ (.D(_0265_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8789_ (.D(_0266_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8790_ (.D(_0267_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8791_ (.D(_0268_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8792_ (.D(_0269_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8793_ (.D(_0270_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8794_ (.D(_0271_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8795_ (.D(_0272_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8796_ (.D(_0273_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8797_ (.D(_0274_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8798_ (.D(_0275_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8799_ (.D(_0276_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8800_ (.D(_0277_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8801_ (.D(_0278_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8802_ (.D(_0279_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8803_ (.D(_0280_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8804_ (.D(_0281_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8805_ (.D(_0282_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8806_ (.D(_0283_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_94 (.Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_89 (.Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8848_ (.I(net46),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8849_ (.I(net46),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8850_ (.I(net46),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8851_ (.I(net46),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8852_ (.I(net47),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8853_ (.I(net47),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8854_ (.I(net47),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[5]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(io_in[6]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input7 (.I(io_in[7]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(io_in[8]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(io_in[9]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(wb_rst_i),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net50),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net53),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net52),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net13),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net36),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net33),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout53 (.I(net29),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_opt_2_1_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_1_wb_clk_i (.I(clknet_opt_2_0_wb_clk_i),
    .Z(clknet_opt_2_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__D (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__D (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__D (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__D (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__D (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__D (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__D (.I(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__D (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__D (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__D (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__D (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__D (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__D (.I(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__D (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__D (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__D (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8725__D (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__D (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__D (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__D (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__D (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__D (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8801__D (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__I (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__S (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__S (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__S1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__S1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A4 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__I (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__B2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__C2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__I (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__I (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__I (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__I (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__B1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A3 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__B1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__C (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__B1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__B1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__A3 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__C (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A3 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__I0 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__B (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__C (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__B2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__C (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__B2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__B2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__B2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__B2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__B (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A4 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__B (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__B (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__B (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I0 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A3 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__B1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__S (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__S (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__S (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__S (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__I (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A3 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__I (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__I (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A2 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__B2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__I (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__B1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__B1 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A3 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A3 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A4 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__B1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__I (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__I (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A3 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__I0 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__I (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__B2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__C2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__B2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__B2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__B (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__C (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__I0 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__B (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__B (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__B2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A2 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__I (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A3 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__B (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__I (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__B1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__I0 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__B (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A4 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A4 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__B1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__B1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__C2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__B1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__B1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__C (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__B (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__I (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__B2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__B2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__B1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__B1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__I (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A3 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A3 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__I (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A3 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__B2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A3 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__B1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__B1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__B1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__B (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__B2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__I (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A3 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__B2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__B2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A1 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__B1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__B1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__B1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__B (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__I0 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A2 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__C (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__S (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__I0 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__B2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A3 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A3 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__B1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A3 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A3 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__B1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__B2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__B (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__B2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__B (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__I (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__B1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__C1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A3 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__B1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__B (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__B2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__I (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A3 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__B1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__B2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__B2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__I (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__B (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__I (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__B1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__B1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A3 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A3 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__I (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A2 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A2 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__A1 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__B (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__I (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__C (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__B1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__B1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__B1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__I (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A3 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__B2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__I (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A3 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__B (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__B (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__I (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__C (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__I (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A3 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A4 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A3 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A3 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A3 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__I (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__I (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__B2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__C (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__C (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__C (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__I (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__S (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__S (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__C1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__S0 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__S0 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__S0 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__S0 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__S1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__S1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__S1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__B1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__I (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__I (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__I (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__B2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__B2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__B2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__I (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__B2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__B2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__B2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__B2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__B2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I0 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__I (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__B2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__B2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__B2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__B2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__B2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__C (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A1 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__B (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__B2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__B2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S0 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__S0 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__S0 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__B (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__S1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__S1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__S1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__B2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__B (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__B2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__B2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__B2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__B2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__I (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__B2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__B2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__B2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__I1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__I (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__I (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A3 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__I (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__B2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__B1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__B1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__C (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__I (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__I (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__C (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__C (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__C (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__I (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__I (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A4 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__I (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__I (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A1 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A4 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A4 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__I (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__I (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A3 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A3 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__B (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__I (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__I (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A3 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__C (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__I (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A3 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__I (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__B (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__I (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__C (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__I (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__I (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__I (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__I (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A3 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__I (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A3 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__I (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A3 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A3 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__B1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__B2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__I (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__I (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__I (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__I (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__I (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__I (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A1 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__B2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I0 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__B2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I1 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__I (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__I (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__C (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__I (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__B (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__I (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7685__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__I (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__I (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__B (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__I0 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__I1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__I (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__I (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__I0 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__I1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__S (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__S (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__S (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__I (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__I (.I(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__I (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__I (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__I (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A2 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I0 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__I0 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__I (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__I0 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__I (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__I (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__I (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__I (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__B (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__I (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__I (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__B (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__B1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A2 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__I (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__I (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__I (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A3 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__I (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__I (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A3 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__B (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__B (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A3 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A3 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__B (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__I (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__B (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__B (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__I (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__I (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__I (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__I (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__I (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__B2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A3 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A3 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A3 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__I (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__C (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__B (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A3 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A3 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A3 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A3 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__I (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A4 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A3 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A3 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A3 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__B (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__I (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A3 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__B1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__C (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__B (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__C (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__B (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__C (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__B (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__B2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__I (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__I (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__B2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__B (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__B (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A3 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A4 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__C (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__C (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__C (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__C2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__I (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A3 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__B1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A3 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A3 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__B2 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__I (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__B1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__I (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__A3 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A4 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__I (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A4 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__C (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__B (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__B1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__A1 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A3 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__B (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__I (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A4 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A3 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__B1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__C (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__B (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A1 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A1 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__B2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__B (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__C (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A3 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__B (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A3 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__I (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A3 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__C (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__I (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__I (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__I (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__B1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A3 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7683__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A4 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__B1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A3 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__B (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A3 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__B (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A3 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__C (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__I (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__I (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__B (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__B (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__B (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A3 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__B (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__I (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__C (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__B (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__I (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__I (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__I (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__B2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__B (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__C (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__I (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__B (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__C (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__I (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__I (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__I (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__B (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__C (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__B (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A3 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A4 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__C (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__B (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__I (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__B1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__C1 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__I (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__B (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__I (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A2 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__A2 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__I (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__I (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__C (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__B (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__S (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__C (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__C (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__C (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__B (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__I (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__I (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__I (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__I (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__C (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__B2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__C (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__B (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__B1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__B2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__I1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__B2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__I (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A1 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__I (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__I (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__I (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__B2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A3 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__I (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A4 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__B (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__B (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__B1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__B2 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__C (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__B1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__B2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__I (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__C2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__B1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__B1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A3 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__C2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__I0 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__B2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__B (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__C (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__I (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__I (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__I (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__I (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__B2 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__I (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__I (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__I (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__I (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A2 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__B (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A1 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__I (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A2 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A2 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__B2 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__I (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__I (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A3 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__I (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__I (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A3 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__C (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__I (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A3 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__I (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A3 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__I (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__I (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__B (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A3 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A3 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__I (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__B (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__C (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__B1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__B1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A3 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__B1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__I (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__I (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A3 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__C (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__B2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A1 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A2 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__B2 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A3 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__I (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__I (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__I (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__S (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__C (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__I (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__B (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A3 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__I (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__I (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__I (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__C (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__C (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__I (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A3 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__I (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A4 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A3 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__C (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__C (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__C (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__I (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__C (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__C (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__I (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__C (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__C (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__C (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__B1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__B (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__B (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__B (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__B (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__C (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__C (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__C (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A4 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__I (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__B (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__B (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__S (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__S (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__B (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__B (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A3 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A3 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__B (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A4 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__C (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__I (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A3 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__C (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__C (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__I (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__B (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__B (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__C (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__C (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A4 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__B2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__B2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__C (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__C (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__C (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__C (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__C (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__B (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__C (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__B (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__C (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A2 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__B1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__C (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__B1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__B2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__B1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A3 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__B1 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__B (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A2 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A2 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__B2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__I0 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__B (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__B (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__B1 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__B1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__B1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__B1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A2 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__B (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__B (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__B (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A3 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__B (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__C (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__B (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__B2 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__B (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A3 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__B (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__C (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__B (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__B1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__B (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A2 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A3 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A4 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A2 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__I (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__I (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__I (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A3 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A2 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A3 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A4 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A2 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__B (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__I (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__I (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A2 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__I (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__I (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A2 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__B2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A3 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A2 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A3 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__I (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A2 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__C (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A3 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A1 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A1 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__B1 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A3 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__I (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__B (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__A1 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__I (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__I (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__B (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__B (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__B (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A2 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A2 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__A1 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A1 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A3 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A1 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__I (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A2 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__I (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A4 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A3 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A4 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__B (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__I (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__I (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__I (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A2 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A2 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__S (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__I (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__I0 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__B (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__I1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A1 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__B2 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__B2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__B2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__B2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__I (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A2 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A2 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A1 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__C (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__I (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A3 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A2 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A3 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__B (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__B (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A2 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A4 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A4 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A2 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__B2 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A1 (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__C (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__C (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__I (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__B (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__B (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__B (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__B (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__B (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A2 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A2 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__C (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__I (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__I (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__B2 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__C (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__A1 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__B (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A1 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__C (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A2 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__B (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__C (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__I (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__I (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__C (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A3 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A2 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A3 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__I (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__B (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__B (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A3 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__C (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__B (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__B (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__B (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__C (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__B1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__I (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A2 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A2 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A2 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A3 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__B (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__B2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A4 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__I (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A2 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__B (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__I (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__B2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__I (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__C (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__A2 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A3 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A4 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A3 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__A1 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A3 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A2 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A1 (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A4 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A1 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A2 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__B (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__C (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A3 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A2 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A3 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A3 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A3 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__A4 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__A1 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A1 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A2 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A2 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A2 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A2 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__A2 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A2 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__A2 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__B (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__B (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__B (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__C (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__B (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A2 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__C (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__I (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__B2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__C (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__C (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__B (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__B2 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A1 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__C (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A2 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A3 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__I (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__B (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__C (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__B (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__B (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__I (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__I (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__I (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__C (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__C (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__C (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__C (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__B1 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A2 (.I(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__B1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A3 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__C (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__A3 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__A2 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A2 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__I (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__C (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__B (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A1 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A1 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A2 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A2 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A4 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__B (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__B2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__C (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A1 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__I (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__B (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__B (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__I (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__B2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__B2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__B1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__I (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__I (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A2 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A2 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A2 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__I (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__I (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__I (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__I (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__C (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A1 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__B (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__B2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__C (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__I (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__C (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A4 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__B (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__I (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__I (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__I (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__I (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__B (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__B (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A2 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__B (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__B2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__B2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__B2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__B (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__B (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__B2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__A2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__B (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__I1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A4 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__I (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__I (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__S (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__S (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__B2 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A1 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A2 (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__B (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__B2 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__C (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A2 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__B (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A1 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__I1 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__B (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__B1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__I1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__I (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__S (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__S (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__S (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A3 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__I (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A2 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A1 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__A2 (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A1 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__B (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__I1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__I1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__B1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A2 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__S (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__C (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__C (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__C (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__I (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__C (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__C (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A3 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__B1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__B (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7512__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__I (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A3 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A3 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__B (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__B1 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__B2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__C (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__C (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__C (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__B2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__C (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__I (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__I (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__B (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__A2 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__C (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__B (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__C (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__C (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__I (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__I (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__C (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__I (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__B1 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__B2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__B2 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__I (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A1 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__B2 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__B (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A2 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A2 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__B2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__C (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__C (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__A2 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__B1 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__C (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__C (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__B (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__C (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__C (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__C (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__C (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__C (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__I (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A1 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__B (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A2 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A1 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__B (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__B (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__B (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__C (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__C (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__C (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__B (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__B (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A2 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__I (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A1 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A1 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A4 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__B (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__C (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A3 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A1 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__I (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__B1 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__B2 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A2 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__B1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__B (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A1 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A1 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__C (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A3 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__A1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__C (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A2 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A2 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__B2 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__C (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A1 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__A1 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A1 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A2 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__B (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A2 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A3 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__C (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__I (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__I (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__I (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A1 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__B1 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__I (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__A1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__B (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__C (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__C (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__B (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__B (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A3 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__B (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__B (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A3 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A2 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__B1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__B (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A4 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A3 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A3 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A3 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__C (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__I (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__B (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__C (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__I (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__I (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__C (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A1 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__I (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__I (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A2 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__I (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__I (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__B2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__B (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__B (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__I (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__I (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__I (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__B2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__B1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__I (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__B2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__B2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__B2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__B2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__C (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__C (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__C (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__C (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__B2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__B2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__B1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__I (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__B2 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__B1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__A2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__B (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A2 (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__I (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__I (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__I (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__I (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A1 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A1 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A1 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__B2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__B (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A2 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A2 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A2 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__B (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__B1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A2 (.I(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__I (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__I (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__I (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A1 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__B2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__I (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__I (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__A1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A2 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__I (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__I (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__I (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__C (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A1 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__B (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__B (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__B (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__B (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__B (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__B (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__I (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__C (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__A1 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A3 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__C (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__C (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__C (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__I (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__B (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__C (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__B (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A1 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__B2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__B2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__B2 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__B2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__I (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__I (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A2 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__B (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__I (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__A1 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__B (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__I (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A3 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__I (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__B2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A1 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__A1 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__B2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A3 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__C (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__I (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__C (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__C (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A2 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__C2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__B2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__A1 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A1 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A1 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A1 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__B2 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__B2 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__B2 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__B2 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__B1 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__B1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__B1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__C (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__C (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__C (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__B2 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__I (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A1 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A2 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A2 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A2 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A2 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__A1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__B (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__B1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A2 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__C (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__I (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A1 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__B (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__C (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__C (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__C (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__A1 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A1 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A1 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__B (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A1 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__C (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A3 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__B (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__B2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__B2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__B1 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__B1 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__B1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__B2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A2 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__B (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__B (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__C (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__C (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A2 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A2 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A2 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__A2 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__B (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__C (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__B (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A1 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__C (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__B (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__B (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__B (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__C (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__B (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__B (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A3 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A2 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__B (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__B (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A1 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__A1 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A1 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__B1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__B1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__B1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__B1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A2 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__B1 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__B2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__B2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A1 (.I(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A1 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__I (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A1 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__B2 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A1 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__A1 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A2 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A2 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__A2 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__B2 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A2 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__B1 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__B1 (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A2 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A2 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__B (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__C (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A1 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__B (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__A2 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__C (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A2 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__B1 (.I(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A2 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A2 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A2 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__A1 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__A3 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A1 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A2 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A2 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A2 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__A1 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__I (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__B (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A1 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__B1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A2 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__C (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__A1 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__I (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__B2 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A1 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__B1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A2 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__A2 (.I(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__B (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__A3 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__C (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__B (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A3 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__A2 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__A1 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A1 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__I (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A1 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__A1 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A1 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__A1 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__B (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A2 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A2 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A2 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__A2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__B1 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A3 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A1 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A1 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__A1 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__C (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__B1 (.I(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A2 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A2 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__B1 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A1 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__I (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A1 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A2 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__B (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__I (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__C (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A1 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A1 (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__B2 (.I(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A1 (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__C (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__C (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__C (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__B (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__I (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A1 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A1 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A1 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A1 (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A1 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__A2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__B1 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A2 (.I(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__B1 (.I(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__B2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A2 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A1 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__A1 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__B (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__B2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__B2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A3 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__B (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__B1 (.I(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__I (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A2 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__B2 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A2 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__I (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A2 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A2 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A2 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__B1 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A1 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A1 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__B2 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__B2 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A1 (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__A1 (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__C (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__C (.I(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__B (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__B2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__B2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__B2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A1 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__B2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__B2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A1 (.I(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A1 (.I(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A1 (.I(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A1 (.I(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__B (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__B (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__B (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__B (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A1 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__A2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__I (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A1 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__A1 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A1 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7532__A1 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A2 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__A2 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__B1 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A1 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A1 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A1 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A1 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__A1 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A1 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__A1 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__B2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A1 (.I(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A1 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__B1 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A2 (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A2 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A2 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A2 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A2 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A1 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A2 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__B (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__B (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__B (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__B (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__B (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A3 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A1 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__A1 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A4 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A3 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A2 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__A2 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__I (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A2 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__B1 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A2 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A2 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__A1 (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A1 (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A1 (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__B (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__B1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A2 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__B (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__I (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__B1 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__B1 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A3 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A2 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__B (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__A1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__C (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__A2 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__B (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__C1 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A2 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A1 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__B1 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__B2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__C (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__B (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__B2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__B1 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__B2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__B1 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A2 (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A2 (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__B (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__B2 (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__B1 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A1 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__I (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__I (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A1 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A3 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__I (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__A2 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A3 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A2 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7685__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7685__A3 (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A3 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A4 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__C (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__C (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__I (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__I (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__B (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A1 (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__B (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__I (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__B (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__I (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__B2 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__B (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A2 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__S (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__I (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__A2 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__I (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__B1 (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__C (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__I (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__I (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__A1 (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A1 (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__C (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__C (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__B1 (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A1 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__C (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__B (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__B2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__C (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A3 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__B (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A1 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A1 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__C (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__B (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__B1 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A2 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A2 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__C (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__B (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__B1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__C (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__C (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__C (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__B (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__A1 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__C (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A1 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A1 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__B (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A2 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A3 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__B (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__C (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__C (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__B (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__B (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__C (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__B (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__C (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__C (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__B2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__C (.I(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__B (.I(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__C (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A2 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__B2 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__B (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__C (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7806__B (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__B (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__B (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__C (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__C (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__C (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__C (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A1 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__C (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__C (.I(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A2 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A2 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A2 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A2 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A2 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__A1 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A1 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A1 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__B (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__I (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__I (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__I (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__I (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__I (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__A2 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A2 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A2 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__A2 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A2 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A2 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A2 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A2 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A2 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__A2 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__A2 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A2 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__A2 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A1 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__A1 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__B2 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A2 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A3 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__I (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__I (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__I (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__I (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__C (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__I (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A1 (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A2 (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__B2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A1 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__B (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A1 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A1 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__B (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__B (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__I (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__B2 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__B (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A2 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__A1 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__A1 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__I (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__B1 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__A1 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__A1 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__B1 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__B1 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__B (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__B1 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__B2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__B2 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__B (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__C (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A1 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__A1 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A2 (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__B (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__I (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__I (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__A2 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A2 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A2 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__A2 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__I (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__I (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__B2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A1 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A1 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__B2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__B1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__B2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__B2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__B2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__B2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A2 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A2 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A2 (.I(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A2 (.I(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__B1 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A1 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A1 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A2 (.I(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__B1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__A1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__B (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__B1 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__A1 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A3 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__B (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A2 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__C (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__B1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__I (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__I (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A2 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A2 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__A2 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A2 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A2 (.I(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__A2 (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__A2 (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A3 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__A2 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__B1 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__B (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A2 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A2 (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A2 (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A2 (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A1 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__C (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A3 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A2 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__A2 (.I(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__B1 (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A2 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__A2 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A2 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A2 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A2 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__B1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__B1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__B1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__B2 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__A2 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__A2 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__I (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A2 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A2 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A2 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A2 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A2 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__A2 (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A2 (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A3 (.I(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__B (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__B (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A2 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A2 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A2 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A2 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__B (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__B (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__B2 (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__B (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__C (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A2 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A3 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__I (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A3 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A1 (.I(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A2 (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A2 (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A3 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__A2 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A2 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__B (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A1 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A2 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A1 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A3 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__B1 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A2 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__A2 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A1 (.I(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A1 (.I(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A2 (.I(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A1 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A1 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__B (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A2 (.I(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A4 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__B1 (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A2 (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A2 (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A2 (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A3 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A3 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__A1 (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__A2 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__A1 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A3 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A2 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__A1 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A2 (.I(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A2 (.I(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__A2 (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__A2 (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A2 (.I(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A2 (.I(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A2 (.I(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__B1 (.I(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__B (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A4 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A2 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A2 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__B1 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__A2 (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__B (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__B1 (.I(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__B (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A1 (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A1 (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__B2 (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A2 (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__A3 (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__I (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__I (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__I (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__I (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__I (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__I (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__I (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__I (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__A1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__B (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__B (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A2 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__B (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A2 (.I(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A1 (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A1 (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A1 (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A1 (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__A1 (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A1 (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A1 (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A1 (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A2 (.I(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A2 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A2 (.I(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A2 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__A3 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A3 (.I(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__A2 (.I(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A3 (.I(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A2 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__A2 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__C (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__B (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A2 (.I(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__B (.I(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__A1 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__I (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A1 (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A2 (.I(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__C (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__A1 (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A3 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A1 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__B (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A2 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__C (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__C (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A1 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A1 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A4 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A2 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A2 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A1 (.I(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__I (.I(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8454__A2 (.I(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__B2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A1 (.I(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__A2 (.I(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A1 (.I(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__A1 (.I(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__B1 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__I (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A3 (.I(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A2 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__B (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A2 (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__B2 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A2 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A3 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A3 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A3 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__B (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__I (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__B (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__B (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A2 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A4 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A4 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__B2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__B (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A2 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A2 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__S0 (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__S0 (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__I (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__S0 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__I (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__S0 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__S0 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__I (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__C2 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__B (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__I (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__B (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__B (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__I (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A1 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__I (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__S (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__S (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__S (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__I (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__S1 (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__S (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__I (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__S (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__S1 (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__S (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__I (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__S1 (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__S (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__S (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__I (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__S1 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__S (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__I (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__S0 (.I(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__S0 (.I(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A1 (.I(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__I (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A2 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__I (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__B (.I(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__I (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__I (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A3 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__I (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__I (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A2 (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A2 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A1 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A1 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A1 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__I (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__I (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__I (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A1 (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__I (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A3 (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A1 (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A2 (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__I (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A1 (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A2 (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A1 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A1 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A2 (.I(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A2 (.I(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A1 (.I(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A1 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A3 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__I (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A2 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A1 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__I (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__I (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A1 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__I (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A3 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A3 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__B (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A1 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A2 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A3 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A3 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A4 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__I (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A1 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A1 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__I (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__I (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__I (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A4 (.I(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__I (.I(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A1 (.I(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A3 (.I(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__I (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__I (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__I (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A2 (.I(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A1 (.I(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A3 (.I(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__B (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A2 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A1 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A1 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A1 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__I (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A1 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A3 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__I (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A1 (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__I (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__I (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A2 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A2 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A2 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__I (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A3 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A3 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A3 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A1 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A2 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A3 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A2 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__I (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A1 (.I(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A1 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__I (.I(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__A2 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__I (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__I (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A3 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__B2 (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__I (.I(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__B (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__A1 (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__I (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__I (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__I (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__B (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A1 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A1 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A3 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A1 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A1 (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A3 (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A3 (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A2 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__I (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A2 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A1 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A2 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A3 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__B (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__I (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A2 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__I (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A3 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__I (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__I (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__I (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A1 (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A2 (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A3 (.I(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A2 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__S (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__I (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__I (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A2 (.I(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A2 (.I(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A3 (.I(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A1 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__B (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__I (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__B (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A3 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A1 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A2 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__C (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__B (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__I (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__I (.I(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A2 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A2 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__I (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__I (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__B (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A2 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__B2 (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I0 (.I(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I1 (.I(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I2 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A2 (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A2 (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I3 (.I(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__I (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__I (.I(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__B (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__I1 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A2 (.I(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__I (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A2 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__C (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__I1 (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__B (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__B2 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__B (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A1 (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A3 (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A1 (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A1 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__B1 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__B (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A1 (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__B2 (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__B (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I (.I(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__B1 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__A1 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__B (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__I (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__C (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A1 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A1 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__B2 (.I(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A2 (.I(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A2 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A2 (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__I (.I(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__A1 (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A2 (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A1 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A3 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A1 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A1 (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__B2 (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__B (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__B (.I(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A3 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A1 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A1 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__B2 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A2 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A1 (.I(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A3 (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A3 (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__B (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__C (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__I (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A2 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__C (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__A1 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A1 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A2 (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A2 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__I (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__I (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A1 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A1 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A1 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A2 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A2 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__I (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__I (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A2 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__I (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A2 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A2 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__B (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__C (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__C (.I(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__I (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A1 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A1 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A3 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A3 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A2 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A2 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A3 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A2 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A3 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A4 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A3 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A3 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__I (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A2 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__I (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A2 (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__B (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__B (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__B (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__B (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A1 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A1 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A1 (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A1 (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__I (.I(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A2 (.I(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A2 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A2 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A2 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A2 (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A2 (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__I (.I(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__A2 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A2 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A3 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A2 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A2 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__B1 (.I(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__B (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__B2 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__B (.I(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__B1 (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__B (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A1 (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__C (.I(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__B (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__C (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__I (.I(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__C (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__B2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A1 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A2 (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__I (.I(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A2 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A3 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A2 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__I (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A1 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__B2 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A3 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A1 (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A1 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__B (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A1 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A3 (.I(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__C (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__A1 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A1 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A2 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__B (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__I (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__B2 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A3 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A2 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A3 (.I(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A2 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__B2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__B2 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A3 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__I (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A3 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__C (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__B (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__I (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__B2 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__B2 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A3 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A2 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A3 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A2 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__I (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A2 (.I(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__B (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__C (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__I (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__C (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__B (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__I (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A1 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__B (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A1 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__C (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__B (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__I (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A2 (.I(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__C (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A1 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__I (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__C (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__C (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__B (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A2 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__I (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__I (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__B2 (.I(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A2 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__I (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__B (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__B2 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__C (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__C (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__B (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__C (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__I (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__B (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__C (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__B2 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A2 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A2 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A2 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A3 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A3 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A3 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__I (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__B2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__B (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A2 (.I(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A1 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__I (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__C (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__I (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__B (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__A2 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A2 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__I (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__A3 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A3 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A2 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__B1 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__B (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__S (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__C (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A1 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A3 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A2 (.I(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A2 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A2 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__I (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A4 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__B1 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A1 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A2 (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A2 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__B1 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A1 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__I (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__I (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__I (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__I (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A1 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__B (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__I (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A4 (.I(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A1 (.I(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A1 (.I(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A3 (.I(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__I (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A2 (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__I (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__S1 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__I (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__I (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A3 (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A3 (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A3 (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__I (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__C1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A3 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A1 (.I(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A1 (.I(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__I (.I(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__I (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A2 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A1 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A1 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__I (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__I (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__I (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__I (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__I (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__I (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__I (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__I (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__I (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__I (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__B (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__B2 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__I (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__I1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__I (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I0 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__I0 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__I (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I0 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__I1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__I3 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I3 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I3 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__B1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A1 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A2 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__B1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__I1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__B1 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I3 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__B2 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__B2 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__B2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A3 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8788__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__CLK (.I(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8765__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8762__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8752__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8758__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8755__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8801__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__CLK (.I(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__CLK (.I(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__CLK (.I(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__CLK (.I(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__CLK (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_1_wb_clk_i_I (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net89;
 assign io_oeb[13] = net94;
 assign io_oeb[14] = net54;
 assign io_oeb[15] = net55;
 assign io_oeb[16] = net56;
 assign io_oeb[17] = net57;
 assign io_oeb[18] = net58;
 assign io_oeb[19] = net59;
 assign io_oeb[1] = net90;
 assign io_oeb[20] = net60;
 assign io_oeb[21] = net61;
 assign io_oeb[22] = net62;
 assign io_oeb[23] = net63;
 assign io_oeb[24] = net64;
 assign io_oeb[25] = net65;
 assign io_oeb[26] = net66;
 assign io_oeb[27] = net67;
 assign io_oeb[28] = net68;
 assign io_oeb[29] = net69;
 assign io_oeb[2] = net91;
 assign io_oeb[30] = net70;
 assign io_oeb[31] = net71;
 assign io_oeb[32] = net72;
 assign io_oeb[33] = net73;
 assign io_oeb[34] = net74;
 assign io_oeb[35] = net75;
 assign io_oeb[36] = net76;
 assign io_oeb[37] = net77;
 assign io_oeb[3] = net92;
 assign io_oeb[4] = net93;
 assign io_out[0] = net78;
 assign io_out[13] = net83;
 assign io_out[1] = net79;
 assign io_out[2] = net80;
 assign io_out[33] = net84;
 assign io_out[34] = net85;
 assign io_out[35] = net86;
 assign io_out[36] = net87;
 assign io_out[37] = net88;
 assign io_out[3] = net81;
 assign io_out[4] = net82;
endmodule

