// This is the unpowered netlist.
module boot_rom (wb_clk_i,
    bus_out,
    cs_port,
    last_addr,
    ram_end,
    ram_start);
 input wb_clk_i;
 output [7:0] bus_out;
 input [2:0] cs_port;
 input [7:0] last_addr;
 input [15:0] ram_end;
 input [15:0] ram_start;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__I (.I(_370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A1 (.I(_362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__A1 (.I(_375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__I (.I(_384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__I (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__I (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__I (.I(_384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__I (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__I (.I(_034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__I (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__I (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__A1 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__A2 (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__B2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__A2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__I (.I(_370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__I (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__C2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__A1 (.I(_375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__I (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__I (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__I (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__I (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__I (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__A1 (.I(_362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__B1 (.I(_092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__A2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__A3 (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__A3 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__A2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__B1 (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__C2 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__552__I (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__B2 (.I(_362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__C2 (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__559__A2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__A2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__B1 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__C2 (.I(_384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__A1 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__I (.I(_034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__B (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__587__A2 (.I(_092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__A1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__A2 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__595__A1 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__598__I (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__599__A2 (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__A2 (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__603__A2 (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__604__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__604__B (.I(_167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__605__A1 (.I(_034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__614__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__615__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__616__C1 (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__616__C2 (.I(_034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__628__A2 (.I(_375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__629__A1 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__629__B2 (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__633__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__634__A1 (.I(_384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__635__A1 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__635__B1 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__641__A1 (.I(_198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__642__A1 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__645__I (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__647__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__653__B1 (.I(_092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__659__I (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__660__C (.I(_167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__662__B (.I(_092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__663__A1 (.I(_370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__665__A1 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__665__B (.I(_375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__671__I (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__672__B1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__673__A2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__675__B1 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__675__B2 (.I(_362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__679__B2 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__682__A2 (.I(_245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__686__A3 (.I(_164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__689__A4 (.I(_252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__692__A3 (.I(_245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__694__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__696__I (.I(_370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__698__B (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__705__A4 (.I(_267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__708__B2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__709__A2 (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__709__B1 (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__713__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__716__A1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__716__A2 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__717__A1 (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__720__A1 (.I(_271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__732__A3 (.I(_289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__734__A1 (.I(_198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__A1 (.I(_296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__747__A2 (.I(_307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__750__C1 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__751__A1 (.I(_198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__751__A4 (.I(_310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__753__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__756__A2 (.I(_167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__761__A1 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__769__A2 (.I(_327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__770__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(last_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(last_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(ram_end[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(ram_end[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(ram_end[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(ram_end[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(ram_end[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(ram_end[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(ram_end[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(ram_end[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(cs_port[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(ram_end[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(ram_end[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(ram_end[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(ram_end[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(ram_end[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(ram_end[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(ram_end[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(ram_end[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(ram_start[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(ram_start[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(cs_port[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(ram_start[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(ram_start[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(ram_start[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(ram_start[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(ram_start[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(ram_start[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(ram_start[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(ram_start[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(ram_start[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(ram_start[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(cs_port[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(ram_start[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(ram_start[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(ram_start[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(ram_start[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(last_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(last_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(last_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(last_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(last_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(last_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _386_ (.I(net3),
    .ZN(_338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _387_ (.A1(net9),
    .A2(net8),
    .ZN(_339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _388_ (.I(_339_),
    .Z(_340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _389_ (.I(net10),
    .Z(_341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _390_ (.I(net11),
    .Z(_342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _391_ (.A1(_341_),
    .A2(_342_),
    .ZN(_343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _392_ (.I(_343_),
    .Z(_344_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _393_ (.A1(_340_),
    .A2(_344_),
    .Z(_345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _394_ (.I(_345_),
    .Z(_346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _395_ (.I(net5),
    .ZN(_347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _396_ (.I(net4),
    .Z(_348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _397_ (.I(_348_),
    .Z(_349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _398_ (.I(net6),
    .ZN(_350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _399_ (.I(_350_),
    .Z(_351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _400_ (.I(net7),
    .Z(_352_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _401_ (.A1(_347_),
    .A2(_349_),
    .A3(_351_),
    .A4(_352_),
    .ZN(_353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _402_ (.I(_353_),
    .Z(_354_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _403_ (.A1(_338_),
    .A2(_346_),
    .A3(_354_),
    .Z(_355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _404_ (.A1(net1),
    .A2(net2),
    .ZN(_356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _405_ (.I(net6),
    .Z(_357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _406_ (.I(net7),
    .ZN(_358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _407_ (.I(_358_),
    .Z(_359_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _408_ (.A1(net5),
    .A2(net4),
    .Z(_360_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _409_ (.A1(_357_),
    .A2(_359_),
    .A3(_360_),
    .ZN(_361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _410_ (.I(_361_),
    .Z(_362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _411_ (.I(net9),
    .Z(_363_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _412_ (.I(_363_),
    .ZN(_364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _413_ (.I(net8),
    .Z(_365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _414_ (.I(_365_),
    .Z(_366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _415_ (.I(_341_),
    .Z(_367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _416_ (.I(net11),
    .ZN(_368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _417_ (.I(_368_),
    .Z(_369_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _418_ (.A1(_364_),
    .A2(_366_),
    .A3(_367_),
    .A4(_369_),
    .ZN(_370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _419_ (.I(_370_),
    .Z(_371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _420_ (.A1(_362_),
    .A2(_371_),
    .ZN(_372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _421_ (.A1(net5),
    .A2(_348_),
    .ZN(_373_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _422_ (.A1(_357_),
    .A2(_359_),
    .A3(_373_),
    .ZN(_374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _423_ (.I(_374_),
    .Z(_375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _424_ (.I(_365_),
    .ZN(_376_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _425_ (.A1(_363_),
    .A2(_376_),
    .A3(_341_),
    .A4(_368_),
    .ZN(_377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _426_ (.I(_377_),
    .Z(_378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _427_ (.I(_378_),
    .Z(_379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _428_ (.A1(_375_),
    .A2(_379_),
    .ZN(_380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _429_ (.I(net5),
    .Z(_381_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _430_ (.I(_348_),
    .ZN(_382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _431_ (.I(_357_),
    .Z(_383_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _432_ (.A1(_381_),
    .A2(_382_),
    .A3(_383_),
    .A4(_359_),
    .ZN(_384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _433_ (.I(_384_),
    .Z(_385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _434_ (.I(_378_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _435_ (.I(_373_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _436_ (.A1(net6),
    .A2(net7),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _437_ (.I(_002_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _438_ (.A1(_001_),
    .A2(_003_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _439_ (.I(_004_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _440_ (.A1(_341_),
    .A2(_369_),
    .A3(_339_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _441_ (.I(_006_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _442_ (.I(_007_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _443_ (.A1(_385_),
    .A2(_000_),
    .B1(_005_),
    .B2(_008_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _444_ (.A1(_372_),
    .A2(_380_),
    .A3(_009_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _445_ (.I(_347_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _446_ (.I(_349_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _447_ (.I(_350_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _448_ (.I(_352_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _449_ (.A1(_011_),
    .A2(_012_),
    .A3(_013_),
    .A4(_014_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _450_ (.A1(_367_),
    .A2(_369_),
    .A3(_340_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _451_ (.I(_384_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _452_ (.I(net10),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _453_ (.I(_018_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _454_ (.I(_342_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _455_ (.A1(_364_),
    .A2(_366_),
    .A3(_019_),
    .A4(_020_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _456_ (.I(_021_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _457_ (.I(_374_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _458_ (.A1(_017_),
    .A2(_022_),
    .B1(_023_),
    .B2(_007_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _459_ (.A1(_015_),
    .A2(_016_),
    .B(_024_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _460_ (.A1(_355_),
    .A2(_356_),
    .B(_010_),
    .C(_025_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _461_ (.I(_363_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _462_ (.A1(_027_),
    .A2(_376_),
    .A3(_018_),
    .A4(_342_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _463_ (.I(_028_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _464_ (.I(_029_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _465_ (.I(_381_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _466_ (.I(_382_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _467_ (.A1(net6),
    .A2(net7),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _468_ (.A1(_031_),
    .A2(_032_),
    .A3(_033_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _469_ (.I(_034_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _470_ (.A1(_031_),
    .A2(_382_),
    .A3(_002_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _471_ (.I(_036_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _472_ (.I(_037_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _473_ (.I(_007_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _474_ (.A1(_030_),
    .A2(_035_),
    .B1(_038_),
    .B2(_039_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _475_ (.I(_022_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _476_ (.A1(_364_),
    .A2(_365_),
    .A3(_343_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _477_ (.I(_042_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _478_ (.I(_043_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _479_ (.A1(_041_),
    .A2(_044_),
    .B(_038_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _480_ (.A1(_340_),
    .A2(_344_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _481_ (.I(_358_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _482_ (.A1(_381_),
    .A2(_349_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _483_ (.A1(_383_),
    .A2(_047_),
    .A3(_048_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _484_ (.A1(_046_),
    .A2(_049_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _485_ (.I(_050_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _486_ (.A1(net42),
    .A2(_051_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _487_ (.I(_345_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _488_ (.I(_028_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _489_ (.I(_360_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _490_ (.A1(_055_),
    .A2(_003_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _491_ (.A1(_053_),
    .A2(_004_),
    .B1(_054_),
    .B2(_056_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _492_ (.A1(_040_),
    .A2(_045_),
    .A3(_052_),
    .A4(_057_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _493_ (.I(_348_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _494_ (.A1(_031_),
    .A2(_059_),
    .A3(_383_),
    .A4(_047_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _495_ (.A1(_046_),
    .A2(_060_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _496_ (.I(_061_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _497_ (.A1(_013_),
    .A2(_014_),
    .A3(_048_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _498_ (.A1(_046_),
    .A2(_063_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _499_ (.I(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _500_ (.A1(net26),
    .A2(_062_),
    .B1(_065_),
    .B2(net12),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _501_ (.I(_370_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _502_ (.A1(_381_),
    .A2(_382_),
    .A3(_351_),
    .A4(_352_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _503_ (.I(_068_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _504_ (.I(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _505_ (.I(_357_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _506_ (.I(_047_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _507_ (.A1(_012_),
    .A2(_071_),
    .A3(_072_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _508_ (.A1(_345_),
    .A2(_068_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _509_ (.I(_074_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _510_ (.A1(_067_),
    .A2(_070_),
    .B1(_073_),
    .B2(_030_),
    .C1(_075_),
    .C2(net28),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _511_ (.A1(_026_),
    .A2(_058_),
    .A3(_066_),
    .A4(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _512_ (.A1(_375_),
    .A2(_054_),
    .B1(_038_),
    .B2(_371_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _513_ (.A1(_347_),
    .A2(_349_),
    .A3(_002_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _514_ (.I(_079_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _515_ (.I(_080_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _516_ (.A1(_019_),
    .A2(_020_),
    .A3(_340_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _517_ (.I(_082_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _518_ (.A1(_371_),
    .A2(_081_),
    .B1(_083_),
    .B2(_005_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _519_ (.A1(_078_),
    .A2(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _520_ (.I(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _521_ (.I(_004_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _522_ (.A1(_067_),
    .A2(_087_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _523_ (.A1(_087_),
    .A2(_035_),
    .B(_379_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _524_ (.I(_082_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _525_ (.A1(_027_),
    .A2(_376_),
    .A3(_344_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _526_ (.I(_091_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _527_ (.I(_033_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _528_ (.A1(_001_),
    .A2(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _529_ (.I(_094_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _530_ (.A1(_363_),
    .A2(_365_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _531_ (.A1(_367_),
    .A2(_020_),
    .A3(_096_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _532_ (.I(_097_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _533_ (.I(_098_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _534_ (.A1(_351_),
    .A2(_014_),
    .A3(_360_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _535_ (.I(_100_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _536_ (.I(_101_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _537_ (.A1(_362_),
    .A2(_090_),
    .B1(_092_),
    .B2(_095_),
    .C1(_099_),
    .C2(_102_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _538_ (.A1(_089_),
    .A2(_103_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _539_ (.A1(_347_),
    .A2(_059_),
    .A3(_033_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _540_ (.I(_105_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _541_ (.A1(_354_),
    .A2(_056_),
    .A3(_106_),
    .B(_098_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _542_ (.I(_091_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _543_ (.A1(_374_),
    .A2(_361_),
    .A3(_056_),
    .A4(_068_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _544_ (.I(_031_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _545_ (.A1(_110_),
    .A2(_032_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _546_ (.A1(_011_),
    .A2(_059_),
    .A3(_071_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _547_ (.A1(_071_),
    .A2(_111_),
    .B(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _548_ (.A1(_029_),
    .A2(_080_),
    .B1(_108_),
    .B2(_109_),
    .C1(_113_),
    .C2(_043_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _549_ (.A1(_107_),
    .A2(_114_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _550_ (.I(_115_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _551_ (.A1(_086_),
    .A2(_088_),
    .A3(_104_),
    .A4(_116_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _552_ (.I(_082_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _553_ (.A1(_017_),
    .A2(_118_),
    .B1(_095_),
    .B2(_029_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _554_ (.A1(_019_),
    .A2(_342_),
    .A3(_096_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _555_ (.I(_120_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _556_ (.I(_377_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _557_ (.A1(_023_),
    .A2(_098_),
    .B1(_121_),
    .B2(_362_),
    .C1(_122_),
    .C2(_100_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _558_ (.A1(_119_),
    .A2(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _559_ (.A1(_023_),
    .A2(_082_),
    .B1(_105_),
    .B2(_120_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _560_ (.A1(_345_),
    .A2(_080_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _561_ (.A1(_021_),
    .A2(_361_),
    .B1(_122_),
    .B2(_354_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _562_ (.A1(_378_),
    .A2(_069_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _563_ (.A1(_125_),
    .A2(_126_),
    .A3(_127_),
    .A4(_128_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _564_ (.A1(_124_),
    .A2(_129_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _565_ (.I(_346_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _566_ (.A1(_011_),
    .A2(_059_),
    .A3(_383_),
    .A4(_359_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _567_ (.I(_132_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _568_ (.A1(_354_),
    .A2(_068_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _569_ (.A1(_351_),
    .A2(_352_),
    .A3(_001_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _570_ (.I(_135_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _571_ (.A1(_054_),
    .A2(_136_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _572_ (.A1(_131_),
    .A2(_133_),
    .B1(_134_),
    .B2(_030_),
    .C(_137_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _573_ (.A1(_055_),
    .A2(_093_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _574_ (.I(_139_),
    .Z(_140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _575_ (.I(_140_),
    .Z(_141_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _576_ (.A1(_036_),
    .A2(_079_),
    .Z(_142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _577_ (.I(_118_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _578_ (.A1(_141_),
    .A2(_142_),
    .B(_143_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _579_ (.A1(_042_),
    .A2(_120_),
    .Z(_145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _580_ (.A1(_122_),
    .A2(_037_),
    .B1(_097_),
    .B2(_139_),
    .C1(_145_),
    .C2(_384_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _581_ (.I(_146_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _582_ (.A1(_138_),
    .A2(_144_),
    .A3(_147_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _583_ (.A1(_043_),
    .A2(_136_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _584_ (.I(_034_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _585_ (.A1(_150_),
    .A2(_080_),
    .B(_108_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _586_ (.A1(_149_),
    .A2(_151_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _587_ (.A1(_102_),
    .A2(_092_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _588_ (.A1(_152_),
    .A2(_153_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _589_ (.A1(_027_),
    .A2(_366_),
    .A3(_367_),
    .A4(_369_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _590_ (.I(_155_),
    .Z(_156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _591_ (.I(_132_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _592_ (.A1(_135_),
    .A2(_139_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _593_ (.A1(_121_),
    .A2(_157_),
    .B1(_158_),
    .B2(_022_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _594_ (.A1(_060_),
    .A2(_156_),
    .B(_159_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _595_ (.A1(_130_),
    .A2(_148_),
    .A3(_154_),
    .A4(_160_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _596_ (.A1(_077_),
    .A2(_117_),
    .A3(_161_),
    .ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _597_ (.A1(_086_),
    .A2(_088_),
    .A3(_104_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _598_ (.I(_006_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _599_ (.A1(_163_),
    .A2(_106_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _600_ (.A1(_116_),
    .A2(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _601_ (.A1(_001_),
    .A2(_093_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _602_ (.A1(_055_),
    .A2(_003_),
    .A3(_155_),
    .B1(_166_),
    .B2(_046_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _603_ (.A1(_163_),
    .A2(_004_),
    .Z(_168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _604_ (.A1(_039_),
    .A2(_070_),
    .B(_167_),
    .C(_168_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _605_ (.A1(_034_),
    .A2(_121_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _606_ (.A1(_378_),
    .A2(_094_),
    .B1(_098_),
    .B2(_132_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _607_ (.A1(_170_),
    .A2(_171_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _608_ (.I(_353_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _609_ (.A1(_173_),
    .A2(_095_),
    .B(_090_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _610_ (.I(_121_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _611_ (.A1(_005_),
    .A2(_099_),
    .B1(_175_),
    .B2(_173_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _612_ (.A1(_174_),
    .A2(_176_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _613_ (.A1(_172_),
    .A2(_177_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _614_ (.I(net2),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _615_ (.A1(net1),
    .A2(_179_),
    .A3(_355_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _616_ (.A1(_007_),
    .A2(_037_),
    .B1(_142_),
    .B2(_021_),
    .C1(_028_),
    .C2(_034_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _617_ (.A1(_146_),
    .A2(_159_),
    .A3(_180_),
    .A4(_181_),
    .Z(_182_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _618_ (.A1(_169_),
    .A2(_178_),
    .A3(_182_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _619_ (.I(_021_),
    .Z(_184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _620_ (.A1(_027_),
    .A2(_366_),
    .A3(_344_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _621_ (.A1(_055_),
    .A2(_093_),
    .A3(_155_),
    .B1(_185_),
    .B2(_015_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _622_ (.A1(_017_),
    .A2(_184_),
    .B1(_173_),
    .B2(_371_),
    .C(_186_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _623_ (.I(_061_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _624_ (.A1(net43),
    .A2(_051_),
    .B1(_188_),
    .B2(net27),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _625_ (.A1(_187_),
    .A2(_189_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _626_ (.A1(_005_),
    .A2(_175_),
    .B1(_157_),
    .B2(_090_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _627_ (.A1(_022_),
    .A2(_150_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _628_ (.A1(_008_),
    .A2(_375_),
    .B(_192_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _629_ (.A1(_053_),
    .A2(_150_),
    .B1(_101_),
    .B2(_108_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _630_ (.A1(_385_),
    .A2(_163_),
    .B1(_083_),
    .B2(_140_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _631_ (.A1(_191_),
    .A2(_193_),
    .A3(_194_),
    .A4(_195_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _632_ (.A1(_012_),
    .A2(_013_),
    .A3(_014_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _633_ (.A1(_110_),
    .A2(_184_),
    .A3(_197_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _634_ (.A1(_384_),
    .A2(_029_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _635_ (.A1(_053_),
    .A2(_157_),
    .B1(_134_),
    .B2(_054_),
    .C(_199_),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _636_ (.I(_064_),
    .Z(_201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _637_ (.I(_074_),
    .Z(_202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _638_ (.A1(net19),
    .A2(_201_),
    .B1(_202_),
    .B2(net35),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _639_ (.I(_122_),
    .Z(_204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _640_ (.A1(_023_),
    .A2(_204_),
    .B1(_037_),
    .B2(_118_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _641_ (.A1(_198_),
    .A2(_200_),
    .A3(_203_),
    .A4(_205_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _642_ (.A1(_130_),
    .A2(_190_),
    .A3(_196_),
    .A4(_206_),
    .Z(_207_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _643_ (.A1(_162_),
    .A2(_165_),
    .A3(_183_),
    .A4(_207_),
    .Z(_208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _644_ (.I(_208_),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _645_ (.I(_056_),
    .Z(_209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _646_ (.I(_136_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _647_ (.A1(_110_),
    .A2(_032_),
    .A3(_013_),
    .A4(_047_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _648_ (.A1(_063_),
    .A2(_211_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _649_ (.I(_204_),
    .Z(_213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _650_ (.A1(_044_),
    .A2(_209_),
    .B1(_210_),
    .B2(_143_),
    .C1(_212_),
    .C2(_213_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _651_ (.I(_017_),
    .Z(_215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _652_ (.A1(_049_),
    .A2(_166_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _653_ (.A1(_215_),
    .A2(_213_),
    .B1(_092_),
    .B2(_133_),
    .C1(_216_),
    .C2(_044_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _654_ (.A1(_152_),
    .A2(_214_),
    .A3(_217_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _655_ (.I(_181_),
    .Z(_219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _656_ (.I(net1),
    .Z(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _657_ (.A1(_220_),
    .A2(_179_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _658_ (.A1(_355_),
    .A2(_221_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _659_ (.I(_106_),
    .Z(_223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _660_ (.A1(_041_),
    .A2(_223_),
    .B(_192_),
    .C(_167_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _661_ (.A1(_115_),
    .A2(_219_),
    .A3(_222_),
    .A4(_224_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _662_ (.A1(_087_),
    .A2(_223_),
    .B(_092_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _663_ (.A1(_370_),
    .A2(_209_),
    .B1(_157_),
    .B2(_204_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _664_ (.A1(_364_),
    .A2(_019_),
    .A3(_020_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _665_ (.A1(_053_),
    .A2(_228_),
    .B(_375_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _666_ (.A1(_150_),
    .A2(_101_),
    .B(_083_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _667_ (.A1(_226_),
    .A2(_227_),
    .A3(_229_),
    .A4(_230_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _668_ (.A1(_000_),
    .A2(_209_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _669_ (.A1(_146_),
    .A2(_232_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _670_ (.A1(_124_),
    .A2(_177_),
    .A3(_231_),
    .A4(_233_),
    .Z(_234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _671_ (.I(_028_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _672_ (.A1(_385_),
    .A2(_235_),
    .B1(_069_),
    .B2(_008_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _673_ (.A1(_235_),
    .A2(_069_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _674_ (.A1(_081_),
    .A2(_083_),
    .B1(_140_),
    .B2(_204_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _675_ (.A1(_163_),
    .A2(_035_),
    .B1(_043_),
    .B2(_362_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _676_ (.A1(_236_),
    .A2(_237_),
    .A3(_238_),
    .A4(_239_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _677_ (.A1(_025_),
    .A2(_085_),
    .A3(_240_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _678_ (.A1(net13),
    .A2(_062_),
    .B1(_065_),
    .B2(net20),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _679_ (.A1(_016_),
    .A2(_063_),
    .B1(_049_),
    .B2(_156_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _680_ (.A1(_095_),
    .A2(_228_),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _681_ (.A1(_376_),
    .A2(_244_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _682_ (.A1(_243_),
    .A2(_245_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _683_ (.I(_050_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _684_ (.I(_136_),
    .Z(_248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _685_ (.A1(_235_),
    .A2(_248_),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _686_ (.A1(_057_),
    .A2(_249_),
    .A3(_164_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _687_ (.A1(net29),
    .A2(_247_),
    .B1(_202_),
    .B2(net36),
    .C(_250_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _688_ (.A1(_241_),
    .A2(_242_),
    .A3(_246_),
    .A4(_251_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _689_ (.A1(_218_),
    .A2(_225_),
    .A3(_234_),
    .A4(_252_),
    .Z(_253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _690_ (.I(_253_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _691_ (.A1(_147_),
    .A2(_219_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _692_ (.A1(_172_),
    .A2(_186_),
    .A3(_245_),
    .Z(_255_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _693_ (.A1(_154_),
    .A2(_254_),
    .A3(_255_),
    .Z(_256_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _694_ (.A1(_220_),
    .A2(net2),
    .A3(_355_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _695_ (.A1(_131_),
    .A2(_223_),
    .B1(_133_),
    .B2(_008_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _696_ (.I(_370_),
    .Z(_259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _697_ (.A1(_259_),
    .A2(_102_),
    .B1(_248_),
    .B2(_000_),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _698_ (.A1(_259_),
    .A2(_379_),
    .B(_070_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _699_ (.A1(_090_),
    .A2(_133_),
    .B1(_197_),
    .B2(_184_),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _700_ (.A1(_258_),
    .A2(_260_),
    .A3(_261_),
    .A4(_262_),
    .Z(_263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _701_ (.A1(_143_),
    .A2(_142_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _702_ (.A1(net30),
    .A2(_051_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _703_ (.A1(_024_),
    .A2(_264_),
    .A3(_230_),
    .A4(_265_),
    .Z(_266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _704_ (.A1(net14),
    .A2(_188_),
    .B1(_202_),
    .B2(net37),
    .C1(_201_),
    .C2(net21),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _705_ (.A1(_257_),
    .A2(_263_),
    .A3(_266_),
    .A4(_267_),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _706_ (.A1(_235_),
    .A2(_101_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _707_ (.A1(_072_),
    .A2(_048_),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _708_ (.A1(_016_),
    .A2(_269_),
    .B1(_270_),
    .B2(_060_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _709_ (.A1(_248_),
    .A2(_108_),
    .B1(_106_),
    .B2(_000_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _710_ (.A1(_081_),
    .A2(_175_),
    .B1(_140_),
    .B2(_044_),
    .ZN(_273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _711_ (.A1(_272_),
    .A2(_273_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _712_ (.A1(_099_),
    .A2(_212_),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _713_ (.A1(_209_),
    .A2(_070_),
    .B(_184_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _714_ (.A1(_275_),
    .A2(_276_),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _715_ (.A1(_125_),
    .A2(_126_),
    .A3(_127_),
    .Z(_278_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _716_ (.A1(_060_),
    .A2(_156_),
    .B(_278_),
    .C(_159_),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _717_ (.A1(_271_),
    .A2(_274_),
    .A3(_277_),
    .A4(_279_),
    .Z(_280_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _718_ (.A1(_165_),
    .A2(_256_),
    .A3(_268_),
    .A4(_280_),
    .Z(_281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _719_ (.I(_281_),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _720_ (.A1(_271_),
    .A2(_274_),
    .A3(_277_),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _721_ (.A1(_144_),
    .A2(_147_),
    .A3(_214_),
    .Z(_283_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _722_ (.A1(_170_),
    .A2(_171_),
    .A3(_227_),
    .Z(_284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _723_ (.A1(_138_),
    .A2(_284_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _724_ (.A1(net31),
    .A2(_051_),
    .B1(_188_),
    .B2(net15),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _725_ (.A1(net22),
    .A2(_201_),
    .B1(_202_),
    .B2(net38),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _726_ (.A1(_259_),
    .A2(_081_),
    .B1(_143_),
    .B2(_087_),
    .C(_243_),
    .ZN(_288_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _727_ (.A1(_187_),
    .A2(_286_),
    .A3(_287_),
    .A4(_288_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _728_ (.A1(net3),
    .A2(_346_),
    .A3(_173_),
    .Z(_290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _729_ (.A1(_356_),
    .A2(_290_),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _730_ (.A1(_385_),
    .A2(_039_),
    .B1(_131_),
    .B2(_035_),
    .C1(_248_),
    .C2(_259_),
    .ZN(_292_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _731_ (.A1(_224_),
    .A2(_291_),
    .A3(_292_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _732_ (.A1(_279_),
    .A2(_285_),
    .A3(_289_),
    .A4(_293_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _733_ (.A1(_116_),
    .A2(_282_),
    .A3(_283_),
    .A4(_294_),
    .ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _734_ (.A1(_198_),
    .A2(_219_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _735_ (.A1(net32),
    .A2(_247_),
    .B1(_188_),
    .B2(net16),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _736_ (.A1(_215_),
    .A2(_141_),
    .B(_131_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _737_ (.A1(_296_),
    .A2(_297_),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _738_ (.A1(_233_),
    .A2(_255_),
    .A3(_295_),
    .A4(_298_),
    .ZN(_299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _739_ (.A1(_030_),
    .A2(_038_),
    .B1(_210_),
    .B2(_379_),
    .ZN(_300_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _740_ (.A1(_016_),
    .A2(_211_),
    .B1(_185_),
    .B2(_112_),
    .C(_300_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _741_ (.A1(_041_),
    .A2(_223_),
    .ZN(_302_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _742_ (.A1(_372_),
    .A2(_153_),
    .A3(_302_),
    .A4(_237_),
    .ZN(_303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _743_ (.A1(_220_),
    .A2(_179_),
    .A3(_290_),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _744_ (.A1(_144_),
    .A2(_159_),
    .A3(_169_),
    .A4(_304_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _745_ (.A1(_215_),
    .A2(_039_),
    .B(_137_),
    .C(_243_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _746_ (.A1(net23),
    .A2(_065_),
    .B1(_075_),
    .B2(net39),
    .ZN(_307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _747_ (.A1(_306_),
    .A2(_307_),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _748_ (.A1(_301_),
    .A2(_303_),
    .A3(_305_),
    .A4(_308_),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _749_ (.A1(_116_),
    .A2(_299_),
    .A3(_309_),
    .ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _750_ (.A1(net17),
    .A2(_062_),
    .B1(_075_),
    .B2(net40),
    .C1(_134_),
    .C2(_067_),
    .ZN(_310_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _751_ (.A1(_198_),
    .A2(_219_),
    .A3(_284_),
    .A4(_310_),
    .Z(_311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _752_ (.A1(_032_),
    .A2(_118_),
    .B(_346_),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _753_ (.A1(_110_),
    .A2(_003_),
    .A3(_312_),
    .Z(_313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _754_ (.A1(_221_),
    .A2(_290_),
    .ZN(_314_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _755_ (.A1(_306_),
    .A2(_313_),
    .A3(_314_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _756_ (.A1(_186_),
    .A2(_167_),
    .ZN(_316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _757_ (.A1(net33),
    .A2(_247_),
    .B1(_201_),
    .B2(net24),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _758_ (.A1(_316_),
    .A2(_317_),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _759_ (.A1(_011_),
    .A2(_012_),
    .A3(_072_),
    .ZN(_319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _760_ (.A1(_102_),
    .A2(_210_),
    .B(_067_),
    .ZN(_320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _761_ (.A1(_156_),
    .A2(_319_),
    .B(_320_),
    .ZN(_321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _762_ (.A1(_213_),
    .A2(_141_),
    .ZN(_322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _763_ (.A1(_213_),
    .A2(_210_),
    .ZN(_323_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _764_ (.A1(_088_),
    .A2(_322_),
    .A3(_244_),
    .A4(_323_),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _765_ (.A1(_315_),
    .A2(_318_),
    .A3(_321_),
    .A4(_324_),
    .ZN(_325_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _766_ (.A1(_283_),
    .A2(_311_),
    .A3(_325_),
    .ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _767_ (.A1(_152_),
    .A2(_200_),
    .A3(_214_),
    .A4(_217_),
    .Z(_326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _768_ (.A1(_071_),
    .A2(_072_),
    .B(_111_),
    .ZN(_327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _769_ (.A1(_041_),
    .A2(_327_),
    .B(_168_),
    .ZN(_328_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _770_ (.A1(_220_),
    .A2(net2),
    .A3(_290_),
    .ZN(_329_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _771_ (.A1(_313_),
    .A2(_329_),
    .Z(_330_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _772_ (.A1(_078_),
    .A2(_147_),
    .A3(_328_),
    .A4(_330_),
    .Z(_331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _773_ (.A1(net18),
    .A2(_062_),
    .B1(_065_),
    .B2(net25),
    .ZN(_332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _774_ (.A1(net34),
    .A2(_247_),
    .B1(_075_),
    .B2(net41),
    .ZN(_333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _775_ (.A1(_332_),
    .A2(_333_),
    .ZN(_334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _776_ (.A1(_215_),
    .A2(_099_),
    .B1(_175_),
    .B2(_141_),
    .ZN(_335_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _777_ (.A1(_040_),
    .A2(_335_),
    .A3(_194_),
    .A4(_205_),
    .ZN(_336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _778_ (.A1(_334_),
    .A2(_336_),
    .ZN(_337_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _779_ (.A1(_282_),
    .A2(_326_),
    .A3(_331_),
    .A4(_337_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(cs_port[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(last_addr[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(last_addr[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(ram_end[0]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(ram_end[10]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(ram_end[11]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(ram_end[12]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(ram_end[13]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(ram_end[14]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(ram_end[15]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(ram_end[1]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(cs_port[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(ram_end[2]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(ram_end[3]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(ram_end[4]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(ram_end[5]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(ram_end[6]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(ram_end[7]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(ram_end[8]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(ram_end[9]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(ram_start[0]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(ram_start[10]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(cs_port[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(ram_start[11]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(ram_start[12]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(ram_start[13]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(ram_start[14]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(ram_start[15]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(ram_start[1]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(ram_start[2]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(ram_start[3]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(ram_start[4]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(ram_start[5]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(last_addr[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(ram_start[6]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(ram_start[7]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(ram_start[8]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(ram_start[9]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(last_addr[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(last_addr[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input7 (.I(last_addr[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(last_addr[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(last_addr[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output44 (.I(net44),
    .Z(bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output45 (.I(net45),
    .Z(bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output46 (.I(net46),
    .Z(bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output47 (.I(net47),
    .Z(bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output48 (.I(net48),
    .Z(bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output49 (.I(net49),
    .Z(bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output50 (.I(net50),
    .Z(bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output51 (.I(net51),
    .Z(bus_out[7]));
endmodule

