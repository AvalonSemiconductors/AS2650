VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sid_top
  CLASS BLOCK ;
  FOREIGN sid_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 750.000 ;
  PIN DAC_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 746.000 17.360 750.000 ;
    END
  END DAC_clk
  PIN DAC_dat_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 746.000 66.640 750.000 ;
    END
  END DAC_dat_1
  PIN DAC_dat_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 746.000 91.280 750.000 ;
    END
  END DAC_dat_2
  PIN DAC_le
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 746.000 42.000 750.000 ;
    END
  END DAC_le
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 746.000 115.920 750.000 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 746.000 140.560 750.000 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 746.000 165.200 750.000 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 189.280 746.000 189.840 750.000 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 746.000 214.480 750.000 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 746.000 239.120 750.000 ;
    END
  END addr[5]
  PIN bus_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 657.440 746.000 658.000 750.000 ;
    END
  END bus_cyc
  PIN bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 746.000 263.760 750.000 ;
    END
  END bus_in[0]
  PIN bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 746.000 288.400 750.000 ;
    END
  END bus_in[1]
  PIN bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 746.000 313.040 750.000 ;
    END
  END bus_in[2]
  PIN bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 746.000 337.680 750.000 ;
    END
  END bus_in[3]
  PIN bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 746.000 362.320 750.000 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 746.000 386.960 750.000 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 411.040 746.000 411.600 750.000 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 746.000 436.240 750.000 ;
    END
  END bus_in[7]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 746.000 460.880 750.000 ;
    END
  END bus_out[0]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 484.960 746.000 485.520 750.000 ;
    END
  END bus_out[1]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 746.000 510.160 750.000 ;
    END
  END bus_out[2]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 746.000 534.800 750.000 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 746.000 559.440 750.000 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 746.000 584.080 750.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 746.000 608.720 750.000 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 632.800 746.000 633.360 750.000 ;
    END
  END bus_out[7]
  PIN bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 746.000 682.640 750.000 ;
    END
  END bus_we
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 746.000 707.280 750.000 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 731.360 746.000 731.920 750.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 733.340 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 733.340 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 733.340 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 743.120 735.690 ;
      LAYER Metal2 ;
        RECT 6.300 745.700 16.500 746.000 ;
        RECT 17.660 745.700 41.140 746.000 ;
        RECT 42.300 745.700 65.780 746.000 ;
        RECT 66.940 745.700 90.420 746.000 ;
        RECT 91.580 745.700 115.060 746.000 ;
        RECT 116.220 745.700 139.700 746.000 ;
        RECT 140.860 745.700 164.340 746.000 ;
        RECT 165.500 745.700 188.980 746.000 ;
        RECT 190.140 745.700 213.620 746.000 ;
        RECT 214.780 745.700 238.260 746.000 ;
        RECT 239.420 745.700 262.900 746.000 ;
        RECT 264.060 745.700 287.540 746.000 ;
        RECT 288.700 745.700 312.180 746.000 ;
        RECT 313.340 745.700 336.820 746.000 ;
        RECT 337.980 745.700 361.460 746.000 ;
        RECT 362.620 745.700 386.100 746.000 ;
        RECT 387.260 745.700 410.740 746.000 ;
        RECT 411.900 745.700 435.380 746.000 ;
        RECT 436.540 745.700 460.020 746.000 ;
        RECT 461.180 745.700 484.660 746.000 ;
        RECT 485.820 745.700 509.300 746.000 ;
        RECT 510.460 745.700 533.940 746.000 ;
        RECT 535.100 745.700 558.580 746.000 ;
        RECT 559.740 745.700 583.220 746.000 ;
        RECT 584.380 745.700 607.860 746.000 ;
        RECT 609.020 745.700 632.500 746.000 ;
        RECT 633.660 745.700 657.140 746.000 ;
        RECT 658.300 745.700 681.780 746.000 ;
        RECT 682.940 745.700 706.420 746.000 ;
        RECT 707.580 745.700 731.060 746.000 ;
        RECT 732.220 745.700 741.860 746.000 ;
        RECT 6.300 15.490 741.860 745.700 ;
      LAYER Metal3 ;
        RECT 6.250 15.540 741.910 733.460 ;
      LAYER Metal4 ;
        RECT 18.060 24.170 21.940 730.150 ;
        RECT 24.140 24.170 98.740 730.150 ;
        RECT 100.940 24.170 175.540 730.150 ;
        RECT 177.740 24.170 252.340 730.150 ;
        RECT 254.540 24.170 329.140 730.150 ;
        RECT 331.340 24.170 405.940 730.150 ;
        RECT 408.140 24.170 482.740 730.150 ;
        RECT 484.940 24.170 559.540 730.150 ;
        RECT 561.740 24.170 636.340 730.150 ;
        RECT 638.540 24.170 713.140 730.150 ;
        RECT 715.340 24.170 721.700 730.150 ;
  END
END sid_top
END LIBRARY

