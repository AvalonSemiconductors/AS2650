magic
tech gf180mcuD
magscale 1 10
timestamp 1700513443
<< nwell >>
rect 1258 50553 53734 51392
rect 1258 50528 17661 50553
rect 1258 49799 31144 49824
rect 1258 48960 53734 49799
rect 1258 47417 53734 48256
rect 1258 47392 10493 47417
rect 1258 46663 13741 46688
rect 1258 45824 53734 46663
rect 1258 45095 26397 45120
rect 1258 44281 53734 45095
rect 1258 44256 7581 44281
rect 1258 42713 53734 43552
rect 1258 42688 15533 42713
rect 1258 41959 27069 41984
rect 1258 41145 53734 41959
rect 1258 41120 8141 41145
rect 1258 40391 22766 40416
rect 1258 39577 53734 40391
rect 1258 39552 6461 39577
rect 1258 38823 12845 38848
rect 1258 38009 53734 38823
rect 1258 37984 33789 38009
rect 1258 37255 2541 37280
rect 1258 36441 53734 37255
rect 1258 36416 47341 36441
rect 1258 35687 36141 35712
rect 1258 34873 53734 35687
rect 1258 34848 2541 34873
rect 1258 34119 21693 34144
rect 1258 33305 53734 34119
rect 1258 33280 26776 33305
rect 1258 32551 2541 32576
rect 1258 31737 53734 32551
rect 1258 31712 10605 31737
rect 1258 30983 16270 31008
rect 1258 30169 53734 30983
rect 1258 30144 2541 30169
rect 1258 29415 14189 29440
rect 1258 28601 53734 29415
rect 1258 28576 32221 28601
rect 1258 27847 2541 27872
rect 1258 27033 53734 27847
rect 1258 27008 14301 27033
rect 1258 26279 28792 26304
rect 1258 25465 53734 26279
rect 1258 25440 31997 25465
rect 1258 24711 2541 24736
rect 1258 23897 53734 24711
rect 1258 23872 14749 23897
rect 1258 23143 52200 23168
rect 1258 22329 53734 23143
rect 1258 22304 2541 22329
rect 1258 21575 14301 21600
rect 1258 20761 53734 21575
rect 1258 20736 10829 20761
rect 1258 20007 18221 20032
rect 1258 19193 53734 20007
rect 1258 19168 2541 19193
rect 1258 18439 6255 18464
rect 1258 17625 53734 18439
rect 1258 17600 18669 17625
rect 1258 16871 2541 16896
rect 1258 16057 53734 16871
rect 1258 16032 10381 16057
rect 1258 15303 19565 15328
rect 1258 14489 53734 15303
rect 1258 14464 40014 14489
rect 1258 13735 2541 13760
rect 1258 12921 53734 13735
rect 1258 12896 31549 12921
rect 1258 12167 51149 12192
rect 1258 11353 53734 12167
rect 1258 11328 2541 11353
rect 1258 10599 20797 10624
rect 1258 9785 53734 10599
rect 1258 9760 4040 9785
rect 1258 9031 45456 9056
rect 1258 8217 53734 9031
rect 1258 8192 8141 8217
rect 1258 7463 6125 7488
rect 1258 6649 53734 7463
rect 1258 6624 14301 6649
rect 1258 5895 34797 5920
rect 1258 5081 53734 5895
rect 1258 5056 9821 5081
rect 1258 4327 20797 4352
rect 1258 3513 53734 4327
rect 1258 3488 25389 3513
<< pwell >>
rect 1258 51392 53734 51830
rect 1258 49824 53734 50528
rect 1258 48256 53734 48960
rect 1258 46688 53734 47392
rect 1258 45120 53734 45824
rect 1258 43552 53734 44256
rect 1258 41984 53734 42688
rect 1258 40416 53734 41120
rect 1258 38848 53734 39552
rect 1258 37280 53734 37984
rect 1258 35712 53734 36416
rect 1258 34144 53734 34848
rect 1258 32576 53734 33280
rect 1258 31008 53734 31712
rect 1258 29440 53734 30144
rect 1258 27872 53734 28576
rect 1258 26304 53734 27008
rect 1258 24736 53734 25440
rect 1258 23168 53734 23872
rect 1258 21600 53734 22304
rect 1258 20032 53734 20736
rect 1258 18464 53734 19168
rect 1258 16896 53734 17600
rect 1258 15328 53734 16032
rect 1258 13760 53734 14464
rect 1258 12192 53734 12896
rect 1258 10624 53734 11328
rect 1258 9056 53734 9760
rect 1258 7488 53734 8192
rect 1258 5920 53734 6624
rect 1258 4352 53734 5056
rect 1258 3050 53734 3488
<< obsm1 >>
rect 1344 3076 53648 51804
<< metal2 >>
rect 13664 54200 13776 55000
rect 41216 54200 41328 55000
rect 2688 0 2800 800
rect 7168 0 7280 800
rect 11648 0 11760 800
rect 16128 0 16240 800
rect 20608 0 20720 800
rect 25088 0 25200 800
rect 29568 0 29680 800
rect 34048 0 34160 800
rect 38528 0 38640 800
rect 43008 0 43120 800
rect 47488 0 47600 800
rect 51968 0 52080 800
<< obsm2 >>
rect 1708 54140 13604 54200
rect 13836 54140 41156 54200
rect 41388 54140 53396 54200
rect 1708 860 53396 54140
rect 1708 800 2628 860
rect 2860 800 7108 860
rect 7340 800 11588 860
rect 11820 800 16068 860
rect 16300 800 20548 860
rect 20780 800 25028 860
rect 25260 800 29508 860
rect 29740 800 33988 860
rect 34220 800 38468 860
rect 38700 800 42948 860
rect 43180 800 47428 860
rect 47660 800 51908 860
rect 52140 800 53396 860
<< metal3 >>
rect 54200 51520 55000 51632
rect 54200 48832 55000 48944
rect 54200 46144 55000 46256
rect 54200 43456 55000 43568
rect 54200 40768 55000 40880
rect 54200 38080 55000 38192
rect 54200 35392 55000 35504
rect 54200 32704 55000 32816
rect 54200 30016 55000 30128
rect 54200 27328 55000 27440
rect 54200 24640 55000 24752
rect 54200 21952 55000 22064
rect 54200 19264 55000 19376
rect 54200 16576 55000 16688
rect 54200 13888 55000 14000
rect 54200 11200 55000 11312
rect 54200 8512 55000 8624
rect 54200 5824 55000 5936
rect 54200 3136 55000 3248
<< obsm3 >>
rect 1698 51692 54200 51772
rect 1698 51460 54140 51692
rect 1698 49004 54200 51460
rect 1698 48772 54140 49004
rect 1698 46316 54200 48772
rect 1698 46084 54140 46316
rect 1698 43628 54200 46084
rect 1698 43396 54140 43628
rect 1698 40940 54200 43396
rect 1698 40708 54140 40940
rect 1698 38252 54200 40708
rect 1698 38020 54140 38252
rect 1698 35564 54200 38020
rect 1698 35332 54140 35564
rect 1698 32876 54200 35332
rect 1698 32644 54140 32876
rect 1698 30188 54200 32644
rect 1698 29956 54140 30188
rect 1698 27500 54200 29956
rect 1698 27268 54140 27500
rect 1698 24812 54200 27268
rect 1698 24580 54140 24812
rect 1698 22124 54200 24580
rect 1698 21892 54140 22124
rect 1698 19436 54200 21892
rect 1698 19204 54140 19436
rect 1698 16748 54200 19204
rect 1698 16516 54140 16748
rect 1698 14060 54200 16516
rect 1698 13828 54140 14060
rect 1698 11372 54200 13828
rect 1698 11140 54140 11372
rect 1698 8684 54200 11140
rect 1698 8452 54140 8684
rect 1698 5996 54200 8452
rect 1698 5764 54140 5996
rect 1698 3308 54200 5764
rect 1698 3108 54140 3308
<< metal4 >>
rect 4448 3076 4768 51804
rect 19808 3076 20128 51804
rect 35168 3076 35488 51804
rect 50528 3076 50848 51804
<< obsm4 >>
rect 21868 3378 35108 50494
rect 35548 3378 46452 50494
<< labels >>
rlabel metal2 s 38528 0 38640 800 6 RXD
port 1 nsew signal input
rlabel metal2 s 34048 0 34160 800 6 TXD
port 2 nsew signal output
rlabel metal3 s 54200 3136 55000 3248 6 addr[0]
port 3 nsew signal input
rlabel metal3 s 54200 5824 55000 5936 6 addr[1]
port 4 nsew signal input
rlabel metal3 s 54200 8512 55000 8624 6 addr[2]
port 5 nsew signal input
rlabel metal2 s 43008 0 43120 800 6 bus_cyc
port 6 nsew signal input
rlabel metal2 s 47488 0 47600 800 6 bus_we
port 7 nsew signal input
rlabel metal3 s 54200 11200 55000 11312 6 data_in[0]
port 8 nsew signal input
rlabel metal3 s 54200 13888 55000 14000 6 data_in[1]
port 9 nsew signal input
rlabel metal3 s 54200 16576 55000 16688 6 data_in[2]
port 10 nsew signal input
rlabel metal3 s 54200 19264 55000 19376 6 data_in[3]
port 11 nsew signal input
rlabel metal3 s 54200 21952 55000 22064 6 data_in[4]
port 12 nsew signal input
rlabel metal3 s 54200 24640 55000 24752 6 data_in[5]
port 13 nsew signal input
rlabel metal3 s 54200 27328 55000 27440 6 data_in[6]
port 14 nsew signal input
rlabel metal3 s 54200 30016 55000 30128 6 data_in[7]
port 15 nsew signal input
rlabel metal3 s 54200 32704 55000 32816 6 data_out[0]
port 16 nsew signal output
rlabel metal3 s 54200 35392 55000 35504 6 data_out[1]
port 17 nsew signal output
rlabel metal3 s 54200 38080 55000 38192 6 data_out[2]
port 18 nsew signal output
rlabel metal3 s 54200 40768 55000 40880 6 data_out[3]
port 19 nsew signal output
rlabel metal3 s 54200 43456 55000 43568 6 data_out[4]
port 20 nsew signal output
rlabel metal3 s 54200 46144 55000 46256 6 data_out[5]
port 21 nsew signal output
rlabel metal3 s 54200 48832 55000 48944 6 data_out[6]
port 22 nsew signal output
rlabel metal3 s 54200 51520 55000 51632 6 data_out[7]
port 23 nsew signal output
rlabel metal2 s 2688 0 2800 800 6 io_in
port 24 nsew signal input
rlabel metal2 s 20608 0 20720 800 6 io_oeb[0]
port 25 nsew signal output
rlabel metal2 s 25088 0 25200 800 6 io_oeb[1]
port 26 nsew signal output
rlabel metal2 s 29568 0 29680 800 6 io_oeb[2]
port 27 nsew signal output
rlabel metal2 s 7168 0 7280 800 6 io_out[0]
port 28 nsew signal output
rlabel metal2 s 11648 0 11760 800 6 io_out[1]
port 29 nsew signal output
rlabel metal2 s 16128 0 16240 800 6 io_out[2]
port 30 nsew signal output
rlabel metal2 s 51968 0 52080 800 6 irq3
port 31 nsew signal output
rlabel metal2 s 41216 54200 41328 55000 6 rst
port 32 nsew signal input
rlabel metal4 s 4448 3076 4768 51804 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 51804 6 vdd
port 33 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 51804 6 vss
port 34 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 51804 6 vss
port 34 nsew ground bidirectional
rlabel metal2 s 13664 54200 13776 55000 6 wb_clk_i
port 35 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 55000 55000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2038696
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/serial_ports/runs/23_11_20_21_48/results/signoff/serial_ports.magic.gds
string GDS_START 283798
<< end >>

